`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/05/08 16:50:57
// Design Name: 
// Module Name: IB_SWU_Addr_Contr_B6
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module IB_SWU_Addr_Contr_B6(
    input                        clk,
    input                        rst_n,
    input    wire     [31:0]     DIN_0, DIN_1, DIN_2,  DIN_3,  DIN_4,  DIN_5,  DIN_6,  DIN_7,
                                 DIN_8, DIN_9, DIN_10, DIN_11, DIN_12, DIN_13, DIN_14, DIN_15,
                                 DIN_16, DIN_17, DIN_18, DIN_19, DIN_20, DIN_21, DIN_22, DIN_23, 
                                 DIN_24, DIN_25, DIN_26, DIN_27, DIN_28, DIN_29, DIN_30, DIN_31,
                                 DIN_32, DIN_33, DIN_34, DIN_35, DIN_36, DIN_37, DIN_38, DIN_39, 
                                 DIN_40, DIN_41, DIN_42, DIN_43, DIN_44, DIN_45, DIN_46, DIN_47, 
                                 DIN_48, DIN_49, DIN_50, DIN_51, DIN_52, DIN_53, DIN_54, DIN_55, 
                                 DIN_56, DIN_57, DIN_58, DIN_59, DIN_60, DIN_61, DIN_62, DIN_63, 
    output   reg      [ 1:0]     ADDR,
    output   reg                 WEA,
    output   reg                 IB_Addr_SWU_work, IB_Addr_SWU_work_Done,
    output   reg      [ 6:0]     Slide_data_0, Slide_data_1, Slide_data_2,  Slide_data_3,  Slide_data_4,  Slide_data_5,  Slide_data_6,  Slide_data_7,
                                 Slide_data_8, Slide_data_9, Slide_data_10, Slide_data_11, Slide_data_12, Slide_data_13, Slide_data_14, Slide_data_15,
                                 Slide_data_16, Slide_data_17, Slide_data_18, Slide_data_19, Slide_data_20, Slide_data_21, Slide_data_22, Slide_data_23, 
                                 Slide_data_24, Slide_data_25, Slide_data_26, Slide_data_27, Slide_data_28, Slide_data_29, Slide_data_30, Slide_data_31,
                                 Slide_data_32, Slide_data_33, Slide_data_34, Slide_data_35, Slide_data_36, Slide_data_37, Slide_data_38, Slide_data_39, 
                                 Slide_data_40, Slide_data_41, Slide_data_42, Slide_data_43, Slide_data_44, Slide_data_45, Slide_data_46, Slide_data_47, 
                                 Slide_data_48, Slide_data_49, Slide_data_50, Slide_data_51, Slide_data_52, Slide_data_53, Slide_data_54, Slide_data_55, 
                                 Slide_data_56, Slide_data_57, Slide_data_58, Slide_data_59, Slide_data_60, Slide_data_61, Slide_data_62, Slide_data_63, 
    output   reg                 PE_EN  //产生第一个7bit的PE阵列输入数据时，代表了PE有效 
);
//*****************************************************基本照搬Block5的SWU代码*****************************************************
reg   [5:0]     cnt;  //
reg   [4:0]     ADDR_d1, ADDR_d2;
//*********由于要padding5，经过测算，ADDR_cnt第一次计数要从0计数到35，以后只需从0计数到25，故用状态机实现*********
reg    [1:0]    current_state, next_state;
parameter       start         = 2'b00,
                cnt_state_1   = 2'b01,
                cnt_state_2   = 2'b10,
                cnt_done      = 2'b11; 

parameter       CNT_1=6'd32, CNT_2=6'd31;
always@(posedge clk or negedge rst_n)begin
    if(!rst_n)
        current_state <= start;
    else
        current_state <= next_state;
end
always@(*)begin
    case(current_state)
        start:begin
                next_state = cnt_state_1;
        end
        cnt_state_1:begin
            if(cnt == CNT_1)begin
                next_state = cnt_state_2;
            end
            else begin 
                next_state = cnt_state_1;
            end
        end
        cnt_state_2:begin
            if(!(ADDR_d2==1 && cnt==28))begin//20是因为Block5的地址4仅有15个有效数据，另外考虑5个padding  block5则是有23个有效数据
                if(cnt == CNT_2)begin
                    next_state = cnt_state_2;
                end
                else begin 
                    next_state = cnt_state_2;
                end
            end else begin
                next_state = cnt_done;
            end
        end
        default: next_state = cnt_done;     
    endcase
end

always@(posedge clk)begin
    case(current_state)
        start:begin
            cnt <= 0;
        end
        cnt_state_1:begin
            if(cnt == CNT_1)begin
                cnt <= 0;
            end
            else begin 
                cnt <= cnt + 1;
            end
        end
        cnt_state_2:begin
            if(cnt == CNT_2)begin
                cnt <= 0;
            end
            else begin 
                cnt <= cnt + 1;
            end
        end
        cnt_done:begin
            cnt <= 0;
        end
        default: cnt <= 0;     
    endcase
end

reg     IB_Addr_SWU_workd1, IB_Addr_SWU_workd2, IB_Addr_SWU_workd3;


always@(posedge clk or negedge rst_n)begin
    if(!rst_n)begin
        IB_Addr_SWU_work <= 0;
        IB_Addr_SWU_work_Done <= 0;
        PE_EN <= 0;
    end
    else begin
        if(ADDR == 0 && cnt == 0)begin
            IB_Addr_SWU_work <= 1;
//            PE_EN <= 1;
        end
        if(ADDR == 0 && cnt == 2)begin
//            IB_Addr_SWU_work <= 1;
            PE_EN <= 1;
        end
        if(ADDR == 1 && cnt == 28)begin
            IB_Addr_SWU_work <= 0;
            IB_Addr_SWU_work_Done <= 1;
        end
    end
end

always@(posedge clk or negedge rst_n)begin
    if(!rst_n)begin
        ADDR <= 0;
    end
    else begin
        if(ADDR ==0 && cnt == (CNT_1-2))begin
            ADDR <= ADDR + 1;
        end
        else begin
            if(ADDR != 0)begin
                if(cnt == 29)begin
                    ADDR <= ADDR + 1;
                end
             end
        end
    end
end

always@(posedge clk)begin
    ADDR_d1 <= ADDR;
    ADDR_d2 <= ADDR_d1;
end

always@(posedge clk or negedge rst_n)begin
    if(!rst_n)begin
        WEA <= 1;
    end
    else begin
        if(!(ADDR_d2==1 && cnt == 28))begin
            if(cnt == 0 && ADDR == 0)begin
                WEA <= 0;
            end
            else if(ADDR==0 && (cnt == CNT_1-2))begin
                WEA <= 0;
            end
            else if(cnt == 29 && ADDR!=0)begin
                WEA <= 0;
            end
            else begin
                WEA <= 1;
            end
        end else begin
            WEA = 1;
        end
    end
end


reg   [ 4:0]     padding_data;
reg   [36:0]     Pad_and_ADDR1_Temp_0, Pad_and_ADDR1_Temp_1, Pad_and_ADDR1_Temp_2, Pad_and_ADDR1_Temp_3, Pad_and_ADDR1_Temp_4, Pad_and_ADDR1_Temp_5, Pad_and_ADDR1_Temp_6, Pad_and_ADDR1_Temp_7, 
                 Pad_and_ADDR1_Temp_8, Pad_and_ADDR1_Temp_9, Pad_and_ADDR1_Temp_10, Pad_and_ADDR1_Temp_11, Pad_and_ADDR1_Temp_12, Pad_and_ADDR1_Temp_13, Pad_and_ADDR1_Temp_14, Pad_and_ADDR1_Temp_15, 
                 Pad_and_ADDR1_Temp_16, Pad_and_ADDR1_Temp_17, Pad_and_ADDR1_Temp_18, Pad_and_ADDR1_Temp_19, Pad_and_ADDR1_Temp_20, Pad_and_ADDR1_Temp_21, Pad_and_ADDR1_Temp_22, Pad_and_ADDR1_Temp_23, 
                 Pad_and_ADDR1_Temp_24, Pad_and_ADDR1_Temp_25, Pad_and_ADDR1_Temp_26, Pad_and_ADDR1_Temp_27, Pad_and_ADDR1_Temp_28, Pad_and_ADDR1_Temp_29, Pad_and_ADDR1_Temp_30, Pad_and_ADDR1_Temp_31,
                 Pad_and_ADDR1_Temp_32, Pad_and_ADDR1_Temp_33, Pad_and_ADDR1_Temp_34, Pad_and_ADDR1_Temp_35, Pad_and_ADDR1_Temp_36, Pad_and_ADDR1_Temp_37, Pad_and_ADDR1_Temp_38, Pad_and_ADDR1_Temp_39, 
                 Pad_and_ADDR1_Temp_40, Pad_and_ADDR1_Temp_41, Pad_and_ADDR1_Temp_42, Pad_and_ADDR1_Temp_43, Pad_and_ADDR1_Temp_44, Pad_and_ADDR1_Temp_45, Pad_and_ADDR1_Temp_46, Pad_and_ADDR1_Temp_47, 
                 Pad_and_ADDR1_Temp_48, Pad_and_ADDR1_Temp_49, Pad_and_ADDR1_Temp_50, Pad_and_ADDR1_Temp_51, Pad_and_ADDR1_Temp_52, Pad_and_ADDR1_Temp_53, Pad_and_ADDR1_Temp_54, Pad_and_ADDR1_Temp_55, 
                 Pad_and_ADDR1_Temp_56, Pad_and_ADDR1_Temp_57, Pad_and_ADDR1_Temp_58, Pad_and_ADDR1_Temp_59, Pad_and_ADDR1_Temp_60, Pad_and_ADDR1_Temp_61, Pad_and_ADDR1_Temp_62, Pad_and_ADDR1_Temp_63;
reg   [ 5:0]     Temp6_0, Temp6_1, Temp6_2, Temp6_3, Temp6_4, Temp6_5, Temp6_6, Temp6_7, Temp6_8, Temp6_9, Temp6_10, Temp6_11, Temp6_12, Temp6_13, Temp6_14, Temp6_15, 
                 Temp6_16, Temp6_17, Temp6_18, Temp6_19, Temp6_20, Temp6_21, Temp6_22, Temp6_23, Temp6_24, Temp6_25, Temp6_26, Temp6_27, Temp6_28, Temp6_29, Temp6_30, Temp6_31,
                 Temp6_32, Temp6_33, Temp6_34, Temp6_35, Temp6_36, Temp6_37, Temp6_38, Temp6_39, Temp6_40, Temp6_41, Temp6_42, Temp6_43, Temp6_44, Temp6_45, Temp6_46, Temp6_47, 
                 Temp6_48, Temp6_49, Temp6_50, Temp6_51, Temp6_52, Temp6_53, Temp6_54, Temp6_55, Temp6_56, Temp6_57, Temp6_58, Temp6_59, Temp6_60, Temp6_61, Temp6_62, Temp6_63;
reg   [37:0]     Temp6_and_Next_ADDR_Data_0, Temp6_and_Next_ADDR_Data_1, Temp6_and_Next_ADDR_Data_2, Temp6_and_Next_ADDR_Data_3, Temp6_and_Next_ADDR_Data_4, Temp6_and_Next_ADDR_Data_5, Temp6_and_Next_ADDR_Data_6, Temp6_and_Next_ADDR_Data_7, 
                 Temp6_and_Next_ADDR_Data_8, Temp6_and_Next_ADDR_Data_9, Temp6_and_Next_ADDR_Data_10, Temp6_and_Next_ADDR_Data_11, Temp6_and_Next_ADDR_Data_12, Temp6_and_Next_ADDR_Data_13, Temp6_and_Next_ADDR_Data_14, Temp6_and_Next_ADDR_Data_15, 
                 Temp6_and_Next_ADDR_Data_16, Temp6_and_Next_ADDR_Data_17, Temp6_and_Next_ADDR_Data_18, Temp6_and_Next_ADDR_Data_19, Temp6_and_Next_ADDR_Data_20, Temp6_and_Next_ADDR_Data_21, Temp6_and_Next_ADDR_Data_22, Temp6_and_Next_ADDR_Data_23, 
                 Temp6_and_Next_ADDR_Data_24, Temp6_and_Next_ADDR_Data_25, Temp6_and_Next_ADDR_Data_26, Temp6_and_Next_ADDR_Data_27, Temp6_and_Next_ADDR_Data_28, Temp6_and_Next_ADDR_Data_29, Temp6_and_Next_ADDR_Data_30, Temp6_and_Next_ADDR_Data_31,
                 Temp6_and_Next_ADDR_Data_32, Temp6_and_Next_ADDR_Data_33, Temp6_and_Next_ADDR_Data_34, Temp6_and_Next_ADDR_Data_35, Temp6_and_Next_ADDR_Data_36, Temp6_and_Next_ADDR_Data_37, Temp6_and_Next_ADDR_Data_38, Temp6_and_Next_ADDR_Data_39, 
                 Temp6_and_Next_ADDR_Data_40, Temp6_and_Next_ADDR_Data_41, Temp6_and_Next_ADDR_Data_42, Temp6_and_Next_ADDR_Data_43, Temp6_and_Next_ADDR_Data_44, Temp6_and_Next_ADDR_Data_45, Temp6_and_Next_ADDR_Data_46, Temp6_and_Next_ADDR_Data_47, 
                 Temp6_and_Next_ADDR_Data_48, Temp6_and_Next_ADDR_Data_49, Temp6_and_Next_ADDR_Data_50, Temp6_and_Next_ADDR_Data_51, Temp6_and_Next_ADDR_Data_52, Temp6_and_Next_ADDR_Data_53, Temp6_and_Next_ADDR_Data_54, Temp6_and_Next_ADDR_Data_55, 
                 Temp6_and_Next_ADDR_Data_56, Temp6_and_Next_ADDR_Data_57, Temp6_and_Next_ADDR_Data_58, Temp6_and_Next_ADDR_Data_59, Temp6_and_Next_ADDR_Data_60, Temp6_and_Next_ADDR_Data_61, Temp6_and_Next_ADDR_Data_62, Temp6_and_Next_ADDR_Data_63;
reg   [10:0]     Temp6_and_five_one_0, Temp6_and_five_one_1, Temp6_and_five_one_2, Temp6_and_five_one_3, Temp6_and_five_one_4, Temp6_and_five_one_5, Temp6_and_five_one_6, Temp6_and_five_one_7, 
                 Temp6_and_five_one_8, Temp6_and_five_one_9, Temp6_and_five_one_10, Temp6_and_five_one_11, Temp6_and_five_one_12, Temp6_and_five_one_13, Temp6_and_five_one_14, Temp6_and_five_one_15, Temp6_and_five_one_16, 
                 Temp6_and_five_one_17, Temp6_and_five_one_18, Temp6_and_five_one_19, Temp6_and_five_one_20, Temp6_and_five_one_21, Temp6_and_five_one_22, Temp6_and_five_one_23, Temp6_and_five_one_24, Temp6_and_five_one_25, 
                 Temp6_and_five_one_26, Temp6_and_five_one_27, Temp6_and_five_one_28, Temp6_and_five_one_29, Temp6_and_five_one_30, Temp6_and_five_one_31, Temp6_and_five_one_32, Temp6_and_five_one_33, Temp6_and_five_one_34, 
                 Temp6_and_five_one_35, Temp6_and_five_one_36, Temp6_and_five_one_37, Temp6_and_five_one_38, Temp6_and_five_one_39, Temp6_and_five_one_40, Temp6_and_five_one_41, Temp6_and_five_one_42, Temp6_and_five_one_43, 
                 Temp6_and_five_one_44, Temp6_and_five_one_45, Temp6_and_five_one_46, Temp6_and_five_one_47, Temp6_and_five_one_48, Temp6_and_five_one_49, Temp6_and_five_one_50, Temp6_and_five_one_51, Temp6_and_five_one_52, 
                 Temp6_and_five_one_53, Temp6_and_five_one_54, Temp6_and_five_one_55, Temp6_and_five_one_56, Temp6_and_five_one_57, Temp6_and_five_one_58, Temp6_and_five_one_59, Temp6_and_five_one_60, Temp6_and_five_one_61, 
                 Temp6_and_five_one_62, Temp6_and_five_one_63;
always@(posedge clk or negedge rst_n)begin
    if(!rst_n)begin
        padding_data <= 5'b11111;
        
        Slide_data_0 <= 0;
        Temp6_0      <= 0;
        Pad_and_ADDR1_Temp_0 <= 0;
        Temp6_and_Next_ADDR_Data_0 <= 0;
        Temp6_and_five_one_0 <= 0;
        
        Slide_data_1 <= 0;
        Temp6_1      <= 0;
        Pad_and_ADDR1_Temp_1 <= 0;
        Temp6_and_Next_ADDR_Data_1 <= 0;
        Temp6_and_five_one_1 <= 0;
        
        Slide_data_2 <= 0;
        Temp6_2      <= 0;
        Pad_and_ADDR1_Temp_2 <= 0;
        Temp6_and_Next_ADDR_Data_2 <= 0;
        Temp6_and_five_one_2 <= 0;
        
        Slide_data_3 <= 0;
        Temp6_3      <= 0;
        Pad_and_ADDR1_Temp_3 <= 0;
        Temp6_and_Next_ADDR_Data_3 <= 0;
        Temp6_and_five_one_3 <= 0;
        
        Slide_data_4 <= 0;
        Temp6_4      <= 0;
        Pad_and_ADDR1_Temp_4 <= 0;
        Temp6_and_Next_ADDR_Data_4 <= 0;
        Temp6_and_five_one_4 <= 0;
        
        Slide_data_5 <= 0;
        Temp6_5      <= 0;
        Pad_and_ADDR1_Temp_5 <= 0;
        Temp6_and_Next_ADDR_Data_5 <= 0;
        Temp6_and_five_one_5 <= 0;
        
        Slide_data_6 <= 0;
        Temp6_6      <= 0;
        Pad_and_ADDR1_Temp_6 <= 0;
        Temp6_and_Next_ADDR_Data_6 <= 0;
        Temp6_and_five_one_6 <= 0;
        
        Slide_data_7 <= 0;
        Temp6_7      <= 0;
        Pad_and_ADDR1_Temp_7 <= 0;
        Temp6_and_Next_ADDR_Data_7 <= 0;
        Temp6_and_five_one_7 <= 0;
        
        Slide_data_8 <= 0;
        Temp6_8      <= 0;
        Pad_and_ADDR1_Temp_8 <= 0;
        Temp6_and_Next_ADDR_Data_8 <= 0;
        Temp6_and_five_one_8 <= 0;
        
        Slide_data_9 <= 0;
        Temp6_9      <= 0;
        Pad_and_ADDR1_Temp_9 <= 0;
        Temp6_and_Next_ADDR_Data_9 <= 0;
        Temp6_and_five_one_9 <= 0;
        
        Slide_data_10 <= 0;
        Temp6_10      <= 0;
        Pad_and_ADDR1_Temp_10 <= 0;
        Temp6_and_Next_ADDR_Data_10 <= 0;
        Temp6_and_five_one_10 <= 0;
        
        Slide_data_11 <= 0;
        Temp6_11      <= 0;
        Pad_and_ADDR1_Temp_11 <= 0;
        Temp6_and_Next_ADDR_Data_11 <= 0;
        Temp6_and_five_one_11 <= 0;
        
        Slide_data_12 <= 0;
        Temp6_12      <= 0;
        Pad_and_ADDR1_Temp_12 <= 0;
        Temp6_and_Next_ADDR_Data_12 <= 0;
        Temp6_and_five_one_12 <= 0;
        
        Slide_data_13 <= 0;
        Temp6_13      <= 0;
        Pad_and_ADDR1_Temp_13 <= 0;
        Temp6_and_Next_ADDR_Data_13 <= 0;
        Temp6_and_five_one_13 <= 0;
        
        Slide_data_14 <= 0;
        Temp6_14      <= 0;
        Pad_and_ADDR1_Temp_14 <= 0;
        Temp6_and_Next_ADDR_Data_14 <= 0;
        Temp6_and_five_one_14 <= 0;
        
        Slide_data_15 <= 0;
        Temp6_15      <= 0;
        Pad_and_ADDR1_Temp_15 <= 0;
        Temp6_and_Next_ADDR_Data_15 <= 0;
        Temp6_and_five_one_15 <= 0;
        
        Slide_data_16 <= 0;
        Temp6_16      <= 0;
        Pad_and_ADDR1_Temp_16 <= 0;
        Temp6_and_Next_ADDR_Data_16 <= 0;
        Temp6_and_five_one_16 <= 0;
        
        Slide_data_17 <= 0;
        Temp6_17      <= 0;
        Pad_and_ADDR1_Temp_17 <= 0;
        Temp6_and_Next_ADDR_Data_17 <= 0;
        Temp6_and_five_one_17 <= 0;
        
        Slide_data_18 <= 0;
        Temp6_18      <= 0;
        Pad_and_ADDR1_Temp_18 <= 0;
        Temp6_and_Next_ADDR_Data_18 <= 0;
        Temp6_and_five_one_18 <= 0;
        
        Slide_data_19 <= 0;
        Temp6_19      <= 0;
        Pad_and_ADDR1_Temp_19 <= 0;
        Temp6_and_Next_ADDR_Data_19 <= 0;
        Temp6_and_five_one_19 <= 0;
        
        Slide_data_20 <= 0;
        Temp6_20      <= 0;
        Pad_and_ADDR1_Temp_20 <= 0;
        Temp6_and_Next_ADDR_Data_20 <= 0;
        Temp6_and_five_one_20 <= 0;
        
        Slide_data_21 <= 0;
        Temp6_21      <= 0;
        Pad_and_ADDR1_Temp_21 <= 0;
        Temp6_and_Next_ADDR_Data_21 <= 0;
        Temp6_and_five_one_21 <= 0;
        
        Slide_data_22 <= 0;
        Temp6_22      <= 0;
        Pad_and_ADDR1_Temp_22 <= 0;
        Temp6_and_Next_ADDR_Data_22 <= 0;
        Temp6_and_five_one_22 <= 0;
        
        Slide_data_23 <= 0;
        Temp6_23      <= 0;
        Pad_and_ADDR1_Temp_23 <= 0;
        Temp6_and_Next_ADDR_Data_23 <= 0;
        Temp6_and_five_one_23 <= 0;
        
        Slide_data_24 <= 0;
        Temp6_24      <= 0;
        Pad_and_ADDR1_Temp_24 <= 0;
        Temp6_and_Next_ADDR_Data_24 <= 0;
        Temp6_and_five_one_24 <= 0;
        
        Slide_data_25 <= 0;
        Temp6_25      <= 0;
        Pad_and_ADDR1_Temp_25 <= 0;
        Temp6_and_Next_ADDR_Data_25 <= 0;
        Temp6_and_five_one_25 <= 0;
        
        Slide_data_26 <= 0;
        Temp6_26      <= 0;
        Pad_and_ADDR1_Temp_26 <= 0;
        Temp6_and_Next_ADDR_Data_26 <= 0;
        Temp6_and_five_one_26 <= 0;
        
        Slide_data_27 <= 0;
        Temp6_27      <= 0;
        Pad_and_ADDR1_Temp_27 <= 0;
        Temp6_and_Next_ADDR_Data_27 <= 0;
        Temp6_and_five_one_27 <= 0;
        
        Slide_data_28 <= 0;
        Temp6_28      <= 0;
        Pad_and_ADDR1_Temp_28 <= 0;
        Temp6_and_Next_ADDR_Data_28 <= 0;
        Temp6_and_five_one_28 <= 0;
        
        Slide_data_29 <= 0;
        Temp6_29      <= 0;
        Pad_and_ADDR1_Temp_29 <= 0;
        Temp6_and_Next_ADDR_Data_29 <= 0;
        Temp6_and_five_one_29 <= 0;
        
        Slide_data_30 <= 0;
        Temp6_30      <= 0;
        Pad_and_ADDR1_Temp_30 <= 0;
        Temp6_and_Next_ADDR_Data_30 <= 0;
        Temp6_and_five_one_30 <= 0;
        
        Slide_data_31 <= 0;
        Temp6_31      <= 0;
        Pad_and_ADDR1_Temp_31 <= 0;
        Temp6_and_Next_ADDR_Data_31 <= 0;
        Temp6_and_five_one_31 <= 0;
        
        Slide_data_32 <= 0;
        Temp6_32      <= 0;
        Pad_and_ADDR1_Temp_32 <= 0;
        Temp6_and_Next_ADDR_Data_32 <= 0;
        Temp6_and_five_one_32 <= 0;
        
        Slide_data_33 <= 0;
        Temp6_33      <= 0;
        Pad_and_ADDR1_Temp_33 <= 0;
        Temp6_and_Next_ADDR_Data_33 <= 0;
        Temp6_and_five_one_33 <= 0;
        
        Slide_data_34 <= 0;
        Temp6_34      <= 0;
        Pad_and_ADDR1_Temp_34 <= 0;
        Temp6_and_Next_ADDR_Data_34 <= 0;
        Temp6_and_five_one_34 <= 0;
        
        Slide_data_35 <= 0;
        Temp6_35      <= 0;
        Pad_and_ADDR1_Temp_35 <= 0;
        Temp6_and_Next_ADDR_Data_35 <= 0;
        Temp6_and_five_one_35 <= 0;
        
        Slide_data_36 <= 0;
        Temp6_36      <= 0;
        Pad_and_ADDR1_Temp_36 <= 0;
        Temp6_and_Next_ADDR_Data_36 <= 0;
        Temp6_and_five_one_36 <= 0;
        
        Slide_data_37 <= 0;
        Temp6_37      <= 0;
        Pad_and_ADDR1_Temp_37 <= 0;
        Temp6_and_Next_ADDR_Data_37 <= 0;
        Temp6_and_five_one_37 <= 0;
        
        Slide_data_38 <= 0;
        Temp6_38      <= 0;
        Pad_and_ADDR1_Temp_38 <= 0;
        Temp6_and_Next_ADDR_Data_38 <= 0;
        Temp6_and_five_one_38 <= 0;
        
        Slide_data_39 <= 0;
        Temp6_39      <= 0;
        Pad_and_ADDR1_Temp_39 <= 0;
        Temp6_and_Next_ADDR_Data_39 <= 0;
        Temp6_and_five_one_39 <= 0;
        
        Slide_data_40 <= 0;
        Temp6_40      <= 0;
        Pad_and_ADDR1_Temp_40 <= 0;
        Temp6_and_Next_ADDR_Data_40 <= 0;
        Temp6_and_five_one_40 <= 0;
        
        Slide_data_41 <= 0;
        Temp6_41      <= 0;
        Pad_and_ADDR1_Temp_41 <= 0;
        Temp6_and_Next_ADDR_Data_41 <= 0;
        Temp6_and_five_one_41 <= 0;
        
        Slide_data_42 <= 0;
        Temp6_42      <= 0;
        Pad_and_ADDR1_Temp_42 <= 0;
        Temp6_and_Next_ADDR_Data_42 <= 0;
        Temp6_and_five_one_42 <= 0;
        
        Slide_data_43 <= 0;
        Temp6_43      <= 0;
        Pad_and_ADDR1_Temp_43 <= 0;
        Temp6_and_Next_ADDR_Data_43 <= 0;
        Temp6_and_five_one_43 <= 0;
        
        Slide_data_44 <= 0;
        Temp6_44      <= 0;
        Pad_and_ADDR1_Temp_44 <= 0;
        Temp6_and_Next_ADDR_Data_44 <= 0;
        Temp6_and_five_one_44 <= 0;
        
        Slide_data_45 <= 0;
        Temp6_45      <= 0;
        Pad_and_ADDR1_Temp_45 <= 0;
        Temp6_and_Next_ADDR_Data_45 <= 0;
        Temp6_and_five_one_45 <= 0;
        
        Slide_data_46 <= 0;
        Temp6_46      <= 0;
        Pad_and_ADDR1_Temp_46 <= 0;
        Temp6_and_Next_ADDR_Data_46 <= 0;
        Temp6_and_five_one_46 <= 0;
        
        Slide_data_47 <= 0;
        Temp6_47      <= 0;
        Pad_and_ADDR1_Temp_47 <= 0;
        Temp6_and_Next_ADDR_Data_47 <= 0;
        Temp6_and_five_one_47 <= 0;
        
        Slide_data_48 <= 0;
        Temp6_48      <= 0;
        Pad_and_ADDR1_Temp_48 <= 0;
        Temp6_and_Next_ADDR_Data_48 <= 0;
        Temp6_and_five_one_48 <= 0;
        
        Slide_data_49 <= 0;
        Temp6_49      <= 0;
        Pad_and_ADDR1_Temp_49 <= 0;
        Temp6_and_Next_ADDR_Data_49 <= 0;
        Temp6_and_five_one_49 <= 0;
        
        Slide_data_50 <= 0;
        Temp6_50      <= 0;
        Pad_and_ADDR1_Temp_50 <= 0;
        Temp6_and_Next_ADDR_Data_50 <= 0;
        Temp6_and_five_one_50 <= 0;
        
        Slide_data_51 <= 0;
        Temp6_51      <= 0;
        Pad_and_ADDR1_Temp_51 <= 0;
        Temp6_and_Next_ADDR_Data_51 <= 0;
        Temp6_and_five_one_51 <= 0;
        
        Slide_data_52 <= 0;
        Temp6_52      <= 0;
        Pad_and_ADDR1_Temp_52 <= 0;
        Temp6_and_Next_ADDR_Data_52 <= 0;
        Temp6_and_five_one_52 <= 0;
        
        Slide_data_53 <= 0;
        Temp6_53      <= 0;
        Pad_and_ADDR1_Temp_53 <= 0;
        Temp6_and_Next_ADDR_Data_53 <= 0;
        Temp6_and_five_one_53 <= 0;
        
        Slide_data_54 <= 0;
        Temp6_54      <= 0;
        Pad_and_ADDR1_Temp_54 <= 0;
        Temp6_and_Next_ADDR_Data_54 <= 0;
        Temp6_and_five_one_54 <= 0;
        
        Slide_data_55 <= 0;
        Temp6_55      <= 0;
        Pad_and_ADDR1_Temp_55 <= 0;
        Temp6_and_Next_ADDR_Data_55 <= 0;
        Temp6_and_five_one_55 <= 0;
        
        Slide_data_56 <= 0;
        Temp6_56      <= 0;
        Pad_and_ADDR1_Temp_56 <= 0;
        Temp6_and_Next_ADDR_Data_56 <= 0;
        Temp6_and_five_one_56 <= 0;
        
        Slide_data_57 <= 0;
        Temp6_57      <= 0;
        Pad_and_ADDR1_Temp_57 <= 0;
        Temp6_and_Next_ADDR_Data_57 <= 0;
        Temp6_and_five_one_57 <= 0;
        
        Slide_data_58 <= 0;
        Temp6_58      <= 0;
        Pad_and_ADDR1_Temp_58 <= 0;
        Temp6_and_Next_ADDR_Data_58 <= 0;
        Temp6_and_five_one_58 <= 0;
        
        Slide_data_59 <= 0;
        Temp6_59      <= 0;
        Pad_and_ADDR1_Temp_59 <= 0;
        Temp6_and_Next_ADDR_Data_59 <= 0;
        Temp6_and_five_one_59 <= 0;
        
        Slide_data_60 <= 0;
        Temp6_60      <= 0;
        Pad_and_ADDR1_Temp_60 <= 0;
        Temp6_and_Next_ADDR_Data_60 <= 0;
        Temp6_and_five_one_60 <= 0;
        
        Slide_data_61 <= 0;
        Temp6_61      <= 0;
        Pad_and_ADDR1_Temp_61 <= 0;
        Temp6_and_Next_ADDR_Data_61 <= 0;
        Temp6_and_five_one_61 <= 0;
        
        Slide_data_62 <= 0;
        Temp6_62      <= 0;
        Pad_and_ADDR1_Temp_62 <= 0;
        Temp6_and_Next_ADDR_Data_62 <= 0;
        Temp6_and_five_one_62 <= 0;
        
        Slide_data_63 <= 0;
        Temp6_63      <= 0;
        Pad_and_ADDR1_Temp_63 <= 0;
        Temp6_and_Next_ADDR_Data_63 <= 0;
        Temp6_and_five_one_63 <= 0;
        

        
    end
    else begin
        if(ADDR_d2 == 0)begin
            if(cnt == 1)begin
                Pad_and_ADDR1_Temp_0 <= {padding_data[4:0], DIN_0[31:0]};
                Temp6_0 <= DIN_0[5:0];
                
                Pad_and_ADDR1_Temp_1 <= {padding_data[4:0], DIN_1[31:0]};
                Temp6_1 <= DIN_1[5:0];
                
                Pad_and_ADDR1_Temp_2 <= {padding_data[4:0], DIN_2[31:0]};
                Temp6_2 <= DIN_2[5:0];
                
                Pad_and_ADDR1_Temp_3 <= {padding_data[4:0], DIN_3[31:0]};
                Temp6_3 <= DIN_3[5:0];
                
                Pad_and_ADDR1_Temp_4 <= {padding_data[4:0], DIN_4[31:0]};
                Temp6_4 <= DIN_4[5:0];
                
                Pad_and_ADDR1_Temp_5 <= {padding_data[4:0], DIN_5[31:0]};
                Temp6_5 <= DIN_5[5:0];
                
                Pad_and_ADDR1_Temp_6 <= {padding_data[4:0], DIN_6[31:0]};
                Temp6_6 <= DIN_6[5:0];
                
                Pad_and_ADDR1_Temp_7 <= {padding_data[4:0], DIN_7[31:0]};
                Temp6_7 <= DIN_7[5:0];
                
                Pad_and_ADDR1_Temp_8 <= {padding_data[4:0], DIN_8[31:0]};
                Temp6_8 <= DIN_8[5:0];
                
                Pad_and_ADDR1_Temp_9 <= {padding_data[4:0], DIN_9[31:0]};
                Temp6_9 <= DIN_9[5:0];
                
                Pad_and_ADDR1_Temp_10 <= {padding_data[4:0], DIN_10[31:0]};
                Temp6_10 <= DIN_10[5:0];
                
                Pad_and_ADDR1_Temp_11 <= {padding_data[4:0], DIN_11[31:0]};
                Temp6_11 <= DIN_11[5:0];
                
                Pad_and_ADDR1_Temp_12 <= {padding_data[4:0], DIN_12[31:0]};
                Temp6_12 <= DIN_12[5:0];
                
                Pad_and_ADDR1_Temp_13 <= {padding_data[4:0], DIN_13[31:0]};
                Temp6_13 <= DIN_13[5:0];
                
                Pad_and_ADDR1_Temp_14 <= {padding_data[4:0], DIN_14[31:0]};
                Temp6_14 <= DIN_14[5:0];
                
                Pad_and_ADDR1_Temp_15 <= {padding_data[4:0], DIN_15[31:0]};
                Temp6_15 <= DIN_15[5:0];
                
                Pad_and_ADDR1_Temp_16 <= {padding_data[4:0], DIN_16[31:0]};
                Temp6_16 <= DIN_16[5:0];
                
                Pad_and_ADDR1_Temp_17 <= {padding_data[4:0], DIN_17[31:0]};
                Temp6_17 <= DIN_17[5:0];
                
                Pad_and_ADDR1_Temp_18 <= {padding_data[4:0], DIN_18[31:0]};
                Temp6_18 <= DIN_18[5:0];
                
                Pad_and_ADDR1_Temp_19 <= {padding_data[4:0], DIN_19[31:0]};
                Temp6_19 <= DIN_19[5:0];
                
                Pad_and_ADDR1_Temp_20 <= {padding_data[4:0], DIN_20[31:0]};
                Temp6_20 <= DIN_20[5:0];
                
                Pad_and_ADDR1_Temp_21 <= {padding_data[4:0], DIN_21[31:0]};
                Temp6_21 <= DIN_21[5:0];
                
                Pad_and_ADDR1_Temp_22 <= {padding_data[4:0], DIN_22[31:0]};
                Temp6_22 <= DIN_22[5:0];
                
                Pad_and_ADDR1_Temp_23 <= {padding_data[4:0], DIN_23[31:0]};
                Temp6_23 <= DIN_23[5:0];
                
                Pad_and_ADDR1_Temp_24 <= {padding_data[4:0], DIN_24[31:0]};
                Temp6_24 <= DIN_24[5:0];
                
                Pad_and_ADDR1_Temp_25 <= {padding_data[4:0], DIN_25[31:0]};
                Temp6_25 <= DIN_25[5:0];
                
                Pad_and_ADDR1_Temp_26 <= {padding_data[4:0], DIN_26[31:0]};
                Temp6_26 <= DIN_26[5:0];
                
                Pad_and_ADDR1_Temp_27 <= {padding_data[4:0], DIN_27[31:0]};
                Temp6_27 <= DIN_27[5:0];
                
                Pad_and_ADDR1_Temp_28 <= {padding_data[4:0], DIN_28[31:0]};
                Temp6_28 <= DIN_28[5:0];
                
                Pad_and_ADDR1_Temp_29 <= {padding_data[4:0], DIN_29[31:0]};
                Temp6_29 <= DIN_29[5:0];
                
                Pad_and_ADDR1_Temp_30 <= {padding_data[4:0], DIN_30[31:0]};
                Temp6_30 <= DIN_30[5:0];
                
                Pad_and_ADDR1_Temp_31 <= {padding_data[4:0], DIN_31[31:0]};
                Temp6_31 <= DIN_31[5:0];
                
                Pad_and_ADDR1_Temp_32 <= {padding_data[4:0], DIN_32[31:0]};
                Temp6_32 <= DIN_32[5:0];
                
                Pad_and_ADDR1_Temp_33 <= {padding_data[4:0], DIN_33[31:0]};
                Temp6_33 <= DIN_33[5:0];
                
                Pad_and_ADDR1_Temp_34 <= {padding_data[4:0], DIN_34[31:0]};
                Temp6_34 <= DIN_34[5:0];
                
                Pad_and_ADDR1_Temp_35 <= {padding_data[4:0], DIN_35[31:0]};
                Temp6_35 <= DIN_35[5:0];
                
                Pad_and_ADDR1_Temp_36 <= {padding_data[4:0], DIN_36[31:0]};
                Temp6_36 <= DIN_36[5:0];
                
                Pad_and_ADDR1_Temp_37 <= {padding_data[4:0], DIN_37[31:0]};
                Temp6_37 <= DIN_37[5:0];
                
                Pad_and_ADDR1_Temp_38 <= {padding_data[4:0], DIN_38[31:0]};
                Temp6_38 <= DIN_38[5:0];
                
                Pad_and_ADDR1_Temp_39 <= {padding_data[4:0], DIN_39[31:0]};
                Temp6_39 <= DIN_39[5:0];
                
                Pad_and_ADDR1_Temp_40 <= {padding_data[4:0], DIN_40[31:0]};
                Temp6_40 <= DIN_40[5:0];
                
                Pad_and_ADDR1_Temp_41 <= {padding_data[4:0], DIN_41[31:0]};
                Temp6_41 <= DIN_41[5:0];
                
                Pad_and_ADDR1_Temp_42 <= {padding_data[4:0], DIN_42[31:0]};
                Temp6_42 <= DIN_42[5:0];
                
                Pad_and_ADDR1_Temp_43 <= {padding_data[4:0], DIN_43[31:0]};
                Temp6_43 <= DIN_43[5:0];
                
                Pad_and_ADDR1_Temp_44 <= {padding_data[4:0], DIN_44[31:0]};
                Temp6_44 <= DIN_44[5:0];
                
                Pad_and_ADDR1_Temp_45 <= {padding_data[4:0], DIN_45[31:0]};
                Temp6_45 <= DIN_45[5:0];
                
                Pad_and_ADDR1_Temp_46 <= {padding_data[4:0], DIN_46[31:0]};
                Temp6_46 <= DIN_46[5:0];
                
                Pad_and_ADDR1_Temp_47 <= {padding_data[4:0], DIN_47[31:0]};
                Temp6_47 <= DIN_47[5:0];
                
                Pad_and_ADDR1_Temp_48 <= {padding_data[4:0], DIN_48[31:0]};
                Temp6_48 <= DIN_48[5:0];
                
                Pad_and_ADDR1_Temp_49 <= {padding_data[4:0], DIN_49[31:0]};
                Temp6_49 <= DIN_49[5:0];
                
                Pad_and_ADDR1_Temp_50 <= {padding_data[4:0], DIN_50[31:0]};
                Temp6_50 <= DIN_50[5:0];
                
                Pad_and_ADDR1_Temp_51 <= {padding_data[4:0], DIN_51[31:0]};
                Temp6_51 <= DIN_51[5:0];
                
                Pad_and_ADDR1_Temp_52 <= {padding_data[4:0], DIN_52[31:0]};
                Temp6_52 <= DIN_52[5:0];
                
                Pad_and_ADDR1_Temp_53 <= {padding_data[4:0], DIN_53[31:0]};
                Temp6_53 <= DIN_53[5:0];
                
                Pad_and_ADDR1_Temp_54 <= {padding_data[4:0], DIN_54[31:0]};
                Temp6_54 <= DIN_54[5:0];
                
                Pad_and_ADDR1_Temp_55 <= {padding_data[4:0], DIN_55[31:0]};
                Temp6_55 <= DIN_55[5:0];
                
                Pad_and_ADDR1_Temp_56 <= {padding_data[4:0], DIN_56[31:0]};
                Temp6_56 <= DIN_56[5:0];
                
                Pad_and_ADDR1_Temp_57 <= {padding_data[4:0], DIN_57[31:0]};
                Temp6_57 <= DIN_57[5:0];
                
                Pad_and_ADDR1_Temp_58 <= {padding_data[4:0], DIN_58[31:0]};
                Temp6_58 <= DIN_58[5:0];
                
                Pad_and_ADDR1_Temp_59 <= {padding_data[4:0], DIN_59[31:0]};
                Temp6_59 <= DIN_59[5:0];
                
                Pad_and_ADDR1_Temp_60 <= {padding_data[4:0], DIN_60[31:0]};
                Temp6_60 <= DIN_60[5:0];
                
                Pad_and_ADDR1_Temp_61 <= {padding_data[4:0], DIN_61[31:0]};
                Temp6_61 <= DIN_61[5:0];
                
                Pad_and_ADDR1_Temp_62 <= {padding_data[4:0], DIN_62[31:0]};
                Temp6_62 <= DIN_62[5:0];
                
                Pad_and_ADDR1_Temp_63 <= {padding_data[4:0], DIN_63[31:0]};
                Temp6_63 <= DIN_63[5:0];            
            end
            else if (cnt <= 32)begin 
                Slide_data_0 <= Pad_and_ADDR1_Temp_0[36:30];
                Pad_and_ADDR1_Temp_0 <= {Pad_and_ADDR1_Temp_0[35:0], 1'b0};
                
                Slide_data_1 <= Pad_and_ADDR1_Temp_1[36:30];
                Pad_and_ADDR1_Temp_1 <= {Pad_and_ADDR1_Temp_1[35:0], 1'b0};
                
                Slide_data_2 <= Pad_and_ADDR1_Temp_2[36:30];
                Pad_and_ADDR1_Temp_2 <= {Pad_and_ADDR1_Temp_2[35:0], 1'b0};
                
                Slide_data_3 <= Pad_and_ADDR1_Temp_3[36:30];
                Pad_and_ADDR1_Temp_3 <= {Pad_and_ADDR1_Temp_3[35:0], 1'b0};
                
                Slide_data_4 <= Pad_and_ADDR1_Temp_4[36:30];
                Pad_and_ADDR1_Temp_4 <= {Pad_and_ADDR1_Temp_4[35:0], 1'b0};
                
                Slide_data_5 <= Pad_and_ADDR1_Temp_5[36:30];
                Pad_and_ADDR1_Temp_5 <= {Pad_and_ADDR1_Temp_5[35:0], 1'b0};
                
                Slide_data_6 <= Pad_and_ADDR1_Temp_6[36:30];
                Pad_and_ADDR1_Temp_6 <= {Pad_and_ADDR1_Temp_6[35:0], 1'b0};
                
                Slide_data_7 <= Pad_and_ADDR1_Temp_7[36:30];
                Pad_and_ADDR1_Temp_7 <= {Pad_and_ADDR1_Temp_7[35:0], 1'b0};
                
                Slide_data_8 <= Pad_and_ADDR1_Temp_8[36:30];
                Pad_and_ADDR1_Temp_8 <= {Pad_and_ADDR1_Temp_8[35:0], 1'b0};
                
                Slide_data_9 <= Pad_and_ADDR1_Temp_9[36:30];
                Pad_and_ADDR1_Temp_9 <= {Pad_and_ADDR1_Temp_9[35:0], 1'b0};
                
                Slide_data_10 <= Pad_and_ADDR1_Temp_10[36:30];
                Pad_and_ADDR1_Temp_10 <= {Pad_and_ADDR1_Temp_10[35:0], 1'b0};
                
                Slide_data_11 <= Pad_and_ADDR1_Temp_11[36:30];
                Pad_and_ADDR1_Temp_11 <= {Pad_and_ADDR1_Temp_11[35:0], 1'b0};
                
                Slide_data_12 <= Pad_and_ADDR1_Temp_12[36:30];
                Pad_and_ADDR1_Temp_12 <= {Pad_and_ADDR1_Temp_12[35:0], 1'b0};
                
                Slide_data_13 <= Pad_and_ADDR1_Temp_13[36:30];
                Pad_and_ADDR1_Temp_13 <= {Pad_and_ADDR1_Temp_13[35:0], 1'b0};
                
                Slide_data_14 <= Pad_and_ADDR1_Temp_14[36:30];
                Pad_and_ADDR1_Temp_14 <= {Pad_and_ADDR1_Temp_14[35:0], 1'b0};
                
                Slide_data_15 <= Pad_and_ADDR1_Temp_15[36:30];
                Pad_and_ADDR1_Temp_15 <= {Pad_and_ADDR1_Temp_15[35:0], 1'b0};
                
                Slide_data_16 <= Pad_and_ADDR1_Temp_16[36:30];
                Pad_and_ADDR1_Temp_16 <= {Pad_and_ADDR1_Temp_16[35:0], 1'b0};
                
                Slide_data_17 <= Pad_and_ADDR1_Temp_17[36:30];
                Pad_and_ADDR1_Temp_17 <= {Pad_and_ADDR1_Temp_17[35:0], 1'b0};
                
                Slide_data_18 <= Pad_and_ADDR1_Temp_18[36:30];
                Pad_and_ADDR1_Temp_18 <= {Pad_and_ADDR1_Temp_18[35:0], 1'b0};
                
                Slide_data_19 <= Pad_and_ADDR1_Temp_19[36:30];
                Pad_and_ADDR1_Temp_19 <= {Pad_and_ADDR1_Temp_19[35:0], 1'b0};
                
                Slide_data_20 <= Pad_and_ADDR1_Temp_20[36:30];
                Pad_and_ADDR1_Temp_20 <= {Pad_and_ADDR1_Temp_20[35:0], 1'b0};
                
                Slide_data_21 <= Pad_and_ADDR1_Temp_21[36:30];
                Pad_and_ADDR1_Temp_21 <= {Pad_and_ADDR1_Temp_21[35:0], 1'b0};
                
                Slide_data_22 <= Pad_and_ADDR1_Temp_22[36:30];
                Pad_and_ADDR1_Temp_22 <= {Pad_and_ADDR1_Temp_22[35:0], 1'b0};
                
                Slide_data_23 <= Pad_and_ADDR1_Temp_23[36:30];
                Pad_and_ADDR1_Temp_23 <= {Pad_and_ADDR1_Temp_23[35:0], 1'b0};
                
                Slide_data_24 <= Pad_and_ADDR1_Temp_24[36:30];
                Pad_and_ADDR1_Temp_24 <= {Pad_and_ADDR1_Temp_24[35:0], 1'b0};
                
                Slide_data_25 <= Pad_and_ADDR1_Temp_25[36:30];
                Pad_and_ADDR1_Temp_25 <= {Pad_and_ADDR1_Temp_25[35:0], 1'b0};
                
                Slide_data_26 <= Pad_and_ADDR1_Temp_26[36:30];
                Pad_and_ADDR1_Temp_26 <= {Pad_and_ADDR1_Temp_26[35:0], 1'b0};
                
                Slide_data_27 <= Pad_and_ADDR1_Temp_27[36:30];
                Pad_and_ADDR1_Temp_27 <= {Pad_and_ADDR1_Temp_27[35:0], 1'b0};
                
                Slide_data_28 <= Pad_and_ADDR1_Temp_28[36:30];
                Pad_and_ADDR1_Temp_28 <= {Pad_and_ADDR1_Temp_28[35:0], 1'b0};
                
                Slide_data_29 <= Pad_and_ADDR1_Temp_29[36:30];
                Pad_and_ADDR1_Temp_29 <= {Pad_and_ADDR1_Temp_29[35:0], 1'b0};
                
                Slide_data_30 <= Pad_and_ADDR1_Temp_30[36:30];
                Pad_and_ADDR1_Temp_30 <= {Pad_and_ADDR1_Temp_30[35:0], 1'b0};
                
                Slide_data_31 <= Pad_and_ADDR1_Temp_31[36:30];
                Pad_and_ADDR1_Temp_31 <= {Pad_and_ADDR1_Temp_31[35:0], 1'b0};
                
                Slide_data_32 <= Pad_and_ADDR1_Temp_32[36:30];
                Pad_and_ADDR1_Temp_32 <= {Pad_and_ADDR1_Temp_32[35:0], 1'b0};
                
                Slide_data_33 <= Pad_and_ADDR1_Temp_33[36:30];
                Pad_and_ADDR1_Temp_33 <= {Pad_and_ADDR1_Temp_33[35:0], 1'b0};
                
                Slide_data_34 <= Pad_and_ADDR1_Temp_34[36:30];
                Pad_and_ADDR1_Temp_34 <= {Pad_and_ADDR1_Temp_34[35:0], 1'b0};
                
                Slide_data_35 <= Pad_and_ADDR1_Temp_35[36:30];
                Pad_and_ADDR1_Temp_35 <= {Pad_and_ADDR1_Temp_35[35:0], 1'b0};
                
                Slide_data_36 <= Pad_and_ADDR1_Temp_36[36:30];
                Pad_and_ADDR1_Temp_36 <= {Pad_and_ADDR1_Temp_36[35:0], 1'b0};
                
                Slide_data_37 <= Pad_and_ADDR1_Temp_37[36:30];
                Pad_and_ADDR1_Temp_37 <= {Pad_and_ADDR1_Temp_37[35:0], 1'b0};
                
                Slide_data_38 <= Pad_and_ADDR1_Temp_38[36:30];
                Pad_and_ADDR1_Temp_38 <= {Pad_and_ADDR1_Temp_38[35:0], 1'b0};
                
                Slide_data_39 <= Pad_and_ADDR1_Temp_39[36:30];
                Pad_and_ADDR1_Temp_39 <= {Pad_and_ADDR1_Temp_39[35:0], 1'b0};
                
                Slide_data_40 <= Pad_and_ADDR1_Temp_40[36:30];
                Pad_and_ADDR1_Temp_40 <= {Pad_and_ADDR1_Temp_40[35:0], 1'b0};
                
                Slide_data_41 <= Pad_and_ADDR1_Temp_41[36:30];
                Pad_and_ADDR1_Temp_41 <= {Pad_and_ADDR1_Temp_41[35:0], 1'b0};
                
                Slide_data_42 <= Pad_and_ADDR1_Temp_42[36:30];
                Pad_and_ADDR1_Temp_42 <= {Pad_and_ADDR1_Temp_42[35:0], 1'b0};
                
                Slide_data_43 <= Pad_and_ADDR1_Temp_43[36:30];
                Pad_and_ADDR1_Temp_43 <= {Pad_and_ADDR1_Temp_43[35:0], 1'b0};
                
                Slide_data_44 <= Pad_and_ADDR1_Temp_44[36:30];
                Pad_and_ADDR1_Temp_44 <= {Pad_and_ADDR1_Temp_44[35:0], 1'b0};
                
                Slide_data_45 <= Pad_and_ADDR1_Temp_45[36:30];
                Pad_and_ADDR1_Temp_45 <= {Pad_and_ADDR1_Temp_45[35:0], 1'b0};
                
                Slide_data_46 <= Pad_and_ADDR1_Temp_46[36:30];
                Pad_and_ADDR1_Temp_46 <= {Pad_and_ADDR1_Temp_46[35:0], 1'b0};
                
                Slide_data_47 <= Pad_and_ADDR1_Temp_47[36:30];
                Pad_and_ADDR1_Temp_47 <= {Pad_and_ADDR1_Temp_47[35:0], 1'b0};
                
                Slide_data_48 <= Pad_and_ADDR1_Temp_48[36:30];
                Pad_and_ADDR1_Temp_48 <= {Pad_and_ADDR1_Temp_48[35:0], 1'b0};
                
                Slide_data_49 <= Pad_and_ADDR1_Temp_49[36:30];
                Pad_and_ADDR1_Temp_49 <= {Pad_and_ADDR1_Temp_49[35:0], 1'b0};
                
                Slide_data_50 <= Pad_and_ADDR1_Temp_50[36:30];
                Pad_and_ADDR1_Temp_50 <= {Pad_and_ADDR1_Temp_50[35:0], 1'b0};
                
                Slide_data_51 <= Pad_and_ADDR1_Temp_51[36:30];
                Pad_and_ADDR1_Temp_51 <= {Pad_and_ADDR1_Temp_51[35:0], 1'b0};
                
                Slide_data_52 <= Pad_and_ADDR1_Temp_52[36:30];
                Pad_and_ADDR1_Temp_52 <= {Pad_and_ADDR1_Temp_52[35:0], 1'b0};
                
                Slide_data_53 <= Pad_and_ADDR1_Temp_53[36:30];
                Pad_and_ADDR1_Temp_53 <= {Pad_and_ADDR1_Temp_53[35:0], 1'b0};
                
                Slide_data_54 <= Pad_and_ADDR1_Temp_54[36:30];
                Pad_and_ADDR1_Temp_54 <= {Pad_and_ADDR1_Temp_54[35:0], 1'b0};
                
                Slide_data_55 <= Pad_and_ADDR1_Temp_55[36:30];
                Pad_and_ADDR1_Temp_55 <= {Pad_and_ADDR1_Temp_55[35:0], 1'b0};
                
                Slide_data_56 <= Pad_and_ADDR1_Temp_56[36:30];
                Pad_and_ADDR1_Temp_56 <= {Pad_and_ADDR1_Temp_56[35:0], 1'b0};
                
                Slide_data_57 <= Pad_and_ADDR1_Temp_57[36:30];
                Pad_and_ADDR1_Temp_57 <= {Pad_and_ADDR1_Temp_57[35:0], 1'b0};
                
                Slide_data_58 <= Pad_and_ADDR1_Temp_58[36:30];
                Pad_and_ADDR1_Temp_58 <= {Pad_and_ADDR1_Temp_58[35:0], 1'b0};
                
                Slide_data_59 <= Pad_and_ADDR1_Temp_59[36:30];
                Pad_and_ADDR1_Temp_59 <= {Pad_and_ADDR1_Temp_59[35:0], 1'b0};
                
                Slide_data_60 <= Pad_and_ADDR1_Temp_60[36:30];
                Pad_and_ADDR1_Temp_60 <= {Pad_and_ADDR1_Temp_60[35:0], 1'b0};
                
                Slide_data_61 <= Pad_and_ADDR1_Temp_61[36:30];
                Pad_and_ADDR1_Temp_61 <= {Pad_and_ADDR1_Temp_61[35:0], 1'b0};
                
                Slide_data_62 <= Pad_and_ADDR1_Temp_62[36:30];
                Pad_and_ADDR1_Temp_62 <= {Pad_and_ADDR1_Temp_62[35:0], 1'b0};
                
                Slide_data_63 <= Pad_and_ADDR1_Temp_63[36:30];
                Pad_and_ADDR1_Temp_63 <= {Pad_and_ADDR1_Temp_63[35:0], 1'b0};              
                if(cnt == 32)begin
                    Temp6_and_Next_ADDR_Data_0 <= {Temp6_0[5:0], DIN_0[31:0]};
                    Temp6_and_Next_ADDR_Data_1 <= {Temp6_1[5:0], DIN_1[31:0]};
                    Temp6_and_Next_ADDR_Data_2 <= {Temp6_2[5:0], DIN_2[31:0]};
                    Temp6_and_Next_ADDR_Data_3 <= {Temp6_3[5:0], DIN_3[31:0]};
                    Temp6_and_Next_ADDR_Data_4 <= {Temp6_4[5:0], DIN_4[31:0]};
                    Temp6_and_Next_ADDR_Data_5 <= {Temp6_5[5:0], DIN_5[31:0]};
                    Temp6_and_Next_ADDR_Data_6 <= {Temp6_6[5:0], DIN_6[31:0]};
                    Temp6_and_Next_ADDR_Data_7 <= {Temp6_7[5:0], DIN_7[31:0]};
                    Temp6_and_Next_ADDR_Data_8 <= {Temp6_8[5:0], DIN_8[31:0]};
                    Temp6_and_Next_ADDR_Data_9 <= {Temp6_9[5:0], DIN_9[31:0]};
                    Temp6_and_Next_ADDR_Data_10 <= {Temp6_10[5:0], DIN_10[31:0]};
                    Temp6_and_Next_ADDR_Data_11 <= {Temp6_11[5:0], DIN_11[31:0]};
                    Temp6_and_Next_ADDR_Data_12 <= {Temp6_12[5:0], DIN_12[31:0]};
                    Temp6_and_Next_ADDR_Data_13 <= {Temp6_13[5:0], DIN_13[31:0]};
                    Temp6_and_Next_ADDR_Data_14 <= {Temp6_14[5:0], DIN_14[31:0]};
                    Temp6_and_Next_ADDR_Data_15 <= {Temp6_15[5:0], DIN_15[31:0]};
                    Temp6_and_Next_ADDR_Data_16 <= {Temp6_16[5:0], DIN_16[31:0]};
                    Temp6_and_Next_ADDR_Data_17 <= {Temp6_17[5:0], DIN_17[31:0]};
                    Temp6_and_Next_ADDR_Data_18 <= {Temp6_18[5:0], DIN_18[31:0]};
                    Temp6_and_Next_ADDR_Data_19 <= {Temp6_19[5:0], DIN_19[31:0]};
                    Temp6_and_Next_ADDR_Data_20 <= {Temp6_20[5:0], DIN_20[31:0]};
                    Temp6_and_Next_ADDR_Data_21 <= {Temp6_21[5:0], DIN_21[31:0]};
                    Temp6_and_Next_ADDR_Data_22 <= {Temp6_22[5:0], DIN_22[31:0]};
                    Temp6_and_Next_ADDR_Data_23 <= {Temp6_23[5:0], DIN_23[31:0]};
                    Temp6_and_Next_ADDR_Data_24 <= {Temp6_24[5:0], DIN_24[31:0]};
                    Temp6_and_Next_ADDR_Data_25 <= {Temp6_25[5:0], DIN_25[31:0]};
                    Temp6_and_Next_ADDR_Data_26 <= {Temp6_26[5:0], DIN_26[31:0]};
                    Temp6_and_Next_ADDR_Data_27 <= {Temp6_27[5:0], DIN_27[31:0]};
                    Temp6_and_Next_ADDR_Data_28 <= {Temp6_28[5:0], DIN_28[31:0]};
                    Temp6_and_Next_ADDR_Data_29 <= {Temp6_29[5:0], DIN_29[31:0]};
                    Temp6_and_Next_ADDR_Data_30 <= {Temp6_30[5:0], DIN_30[31:0]};
                    Temp6_and_Next_ADDR_Data_31 <= {Temp6_31[5:0], DIN_31[31:0]};
                    Temp6_and_Next_ADDR_Data_32 <= {Temp6_32[5:0], DIN_32[31:0]};
                    Temp6_and_Next_ADDR_Data_33 <= {Temp6_33[5:0], DIN_33[31:0]};
                    Temp6_and_Next_ADDR_Data_34 <= {Temp6_34[5:0], DIN_34[31:0]};
                    Temp6_and_Next_ADDR_Data_35 <= {Temp6_35[5:0], DIN_35[31:0]};
                    Temp6_and_Next_ADDR_Data_36 <= {Temp6_36[5:0], DIN_36[31:0]};
                    Temp6_and_Next_ADDR_Data_37 <= {Temp6_37[5:0], DIN_37[31:0]};
                    Temp6_and_Next_ADDR_Data_38 <= {Temp6_38[5:0], DIN_38[31:0]};
                    Temp6_and_Next_ADDR_Data_39 <= {Temp6_39[5:0], DIN_39[31:0]};
                    Temp6_and_Next_ADDR_Data_40 <= {Temp6_40[5:0], DIN_40[31:0]};
                    Temp6_and_Next_ADDR_Data_41 <= {Temp6_41[5:0], DIN_41[31:0]};
                    Temp6_and_Next_ADDR_Data_42 <= {Temp6_42[5:0], DIN_42[31:0]};
                    Temp6_and_Next_ADDR_Data_43 <= {Temp6_43[5:0], DIN_43[31:0]};
                    Temp6_and_Next_ADDR_Data_44 <= {Temp6_44[5:0], DIN_44[31:0]};
                    Temp6_and_Next_ADDR_Data_45 <= {Temp6_45[5:0], DIN_45[31:0]};
                    Temp6_and_Next_ADDR_Data_46 <= {Temp6_46[5:0], DIN_46[31:0]};
                    Temp6_and_Next_ADDR_Data_47 <= {Temp6_47[5:0], DIN_47[31:0]};
                    Temp6_and_Next_ADDR_Data_48 <= {Temp6_48[5:0], DIN_48[31:0]};
                    Temp6_and_Next_ADDR_Data_49 <= {Temp6_49[5:0], DIN_49[31:0]};
                    Temp6_and_Next_ADDR_Data_50 <= {Temp6_50[5:0], DIN_50[31:0]};
                    Temp6_and_Next_ADDR_Data_51 <= {Temp6_51[5:0], DIN_51[31:0]};
                    Temp6_and_Next_ADDR_Data_52 <= {Temp6_52[5:0], DIN_52[31:0]};
                    Temp6_and_Next_ADDR_Data_53 <= {Temp6_53[5:0], DIN_53[31:0]};
                    Temp6_and_Next_ADDR_Data_54 <= {Temp6_54[5:0], DIN_54[31:0]};
                    Temp6_and_Next_ADDR_Data_55 <= {Temp6_55[5:0], DIN_55[31:0]};
                    Temp6_and_Next_ADDR_Data_56 <= {Temp6_56[5:0], DIN_56[31:0]};
                    Temp6_and_Next_ADDR_Data_57 <= {Temp6_57[5:0], DIN_57[31:0]};
                    Temp6_and_Next_ADDR_Data_58 <= {Temp6_58[5:0], DIN_58[31:0]};
                    Temp6_and_Next_ADDR_Data_59 <= {Temp6_59[5:0], DIN_59[31:0]};
                    Temp6_and_Next_ADDR_Data_60 <= {Temp6_60[5:0], DIN_60[31:0]};
                    Temp6_and_Next_ADDR_Data_61 <= {Temp6_61[5:0], DIN_61[31:0]};
                    Temp6_and_Next_ADDR_Data_62 <= {Temp6_62[5:0], DIN_62[31:0]};
                    Temp6_and_Next_ADDR_Data_63 <= {Temp6_63[5:0], DIN_63[31:0]};

                    
                end
             end
         end
         else if(ADDR_d2 == 1)begin
           if(cnt <= 22)begin
                Slide_data_0 <= Temp6_and_Next_ADDR_Data_0[37:31];
                Temp6_and_Next_ADDR_Data_0 <= {Temp6_and_Next_ADDR_Data_0[36:0], 1'b0};
                
                Slide_data_1 <= Temp6_and_Next_ADDR_Data_1[37:31];
                Temp6_and_Next_ADDR_Data_1 <= {Temp6_and_Next_ADDR_Data_1[36:0], 1'b0};
                
                Slide_data_2 <= Temp6_and_Next_ADDR_Data_2[37:31];
                Temp6_and_Next_ADDR_Data_2 <= {Temp6_and_Next_ADDR_Data_2[36:0], 1'b0};
                
                Slide_data_3 <= Temp6_and_Next_ADDR_Data_3[37:31];
                Temp6_and_Next_ADDR_Data_3 <= {Temp6_and_Next_ADDR_Data_3[36:0], 1'b0};
                
                Slide_data_4 <= Temp6_and_Next_ADDR_Data_4[37:31];
                Temp6_and_Next_ADDR_Data_4 <= {Temp6_and_Next_ADDR_Data_4[36:0], 1'b0};
                
                Slide_data_5 <= Temp6_and_Next_ADDR_Data_5[37:31];
                Temp6_and_Next_ADDR_Data_5 <= {Temp6_and_Next_ADDR_Data_5[36:0], 1'b0};
                
                Slide_data_6 <= Temp6_and_Next_ADDR_Data_6[37:31];
                Temp6_and_Next_ADDR_Data_6 <= {Temp6_and_Next_ADDR_Data_6[36:0], 1'b0};
                
                Slide_data_7 <= Temp6_and_Next_ADDR_Data_7[37:31];
                Temp6_and_Next_ADDR_Data_7 <= {Temp6_and_Next_ADDR_Data_7[36:0], 1'b0};
                
                Slide_data_8 <= Temp6_and_Next_ADDR_Data_8[37:31];
                Temp6_and_Next_ADDR_Data_8 <= {Temp6_and_Next_ADDR_Data_8[36:0], 1'b0};
                
                Slide_data_9 <= Temp6_and_Next_ADDR_Data_9[37:31];
                Temp6_and_Next_ADDR_Data_9 <= {Temp6_and_Next_ADDR_Data_9[36:0], 1'b0};
                
                Slide_data_10 <= Temp6_and_Next_ADDR_Data_10[37:31];
                Temp6_and_Next_ADDR_Data_10 <= {Temp6_and_Next_ADDR_Data_10[36:0], 1'b0};
                
                Slide_data_11 <= Temp6_and_Next_ADDR_Data_11[37:31];
                Temp6_and_Next_ADDR_Data_11 <= {Temp6_and_Next_ADDR_Data_11[36:0], 1'b0};
                
                Slide_data_12 <= Temp6_and_Next_ADDR_Data_12[37:31];
                Temp6_and_Next_ADDR_Data_12 <= {Temp6_and_Next_ADDR_Data_12[36:0], 1'b0};
                
                Slide_data_13 <= Temp6_and_Next_ADDR_Data_13[37:31];
                Temp6_and_Next_ADDR_Data_13 <= {Temp6_and_Next_ADDR_Data_13[36:0], 1'b0};
                
                Slide_data_14 <= Temp6_and_Next_ADDR_Data_14[37:31];
                Temp6_and_Next_ADDR_Data_14 <= {Temp6_and_Next_ADDR_Data_14[36:0], 1'b0};
                
                Slide_data_15 <= Temp6_and_Next_ADDR_Data_15[37:31];
                Temp6_and_Next_ADDR_Data_15 <= {Temp6_and_Next_ADDR_Data_15[36:0], 1'b0};
                
                Slide_data_16 <= Temp6_and_Next_ADDR_Data_16[37:31];
                Temp6_and_Next_ADDR_Data_16 <= {Temp6_and_Next_ADDR_Data_16[36:0], 1'b0};
                
                Slide_data_17 <= Temp6_and_Next_ADDR_Data_17[37:31];
                Temp6_and_Next_ADDR_Data_17 <= {Temp6_and_Next_ADDR_Data_17[36:0], 1'b0};
                
                Slide_data_18 <= Temp6_and_Next_ADDR_Data_18[37:31];
                Temp6_and_Next_ADDR_Data_18 <= {Temp6_and_Next_ADDR_Data_18[36:0], 1'b0};
                
                Slide_data_19 <= Temp6_and_Next_ADDR_Data_19[37:31];
                Temp6_and_Next_ADDR_Data_19 <= {Temp6_and_Next_ADDR_Data_19[36:0], 1'b0};
                
                Slide_data_20 <= Temp6_and_Next_ADDR_Data_20[37:31];
                Temp6_and_Next_ADDR_Data_20 <= {Temp6_and_Next_ADDR_Data_20[36:0], 1'b0};
                
                Slide_data_21 <= Temp6_and_Next_ADDR_Data_21[37:31];
                Temp6_and_Next_ADDR_Data_21 <= {Temp6_and_Next_ADDR_Data_21[36:0], 1'b0};
                
                Slide_data_22 <= Temp6_and_Next_ADDR_Data_22[37:31];
                Temp6_and_Next_ADDR_Data_22 <= {Temp6_and_Next_ADDR_Data_22[36:0], 1'b0};
                
                Slide_data_23 <= Temp6_and_Next_ADDR_Data_23[37:31];
                Temp6_and_Next_ADDR_Data_23 <= {Temp6_and_Next_ADDR_Data_23[36:0], 1'b0};
                
                Slide_data_24 <= Temp6_and_Next_ADDR_Data_24[37:31];
                Temp6_and_Next_ADDR_Data_24 <= {Temp6_and_Next_ADDR_Data_24[36:0], 1'b0};
                
                Slide_data_25 <= Temp6_and_Next_ADDR_Data_25[37:31];
                Temp6_and_Next_ADDR_Data_25 <= {Temp6_and_Next_ADDR_Data_25[36:0], 1'b0};
                
                Slide_data_26 <= Temp6_and_Next_ADDR_Data_26[37:31];
                Temp6_and_Next_ADDR_Data_26 <= {Temp6_and_Next_ADDR_Data_26[36:0], 1'b0};
                
                Slide_data_27 <= Temp6_and_Next_ADDR_Data_27[37:31];
                Temp6_and_Next_ADDR_Data_27 <= {Temp6_and_Next_ADDR_Data_27[36:0], 1'b0};
                
                Slide_data_28 <= Temp6_and_Next_ADDR_Data_28[37:31];
                Temp6_and_Next_ADDR_Data_28 <= {Temp6_and_Next_ADDR_Data_28[36:0], 1'b0};
                
                Slide_data_29 <= Temp6_and_Next_ADDR_Data_29[37:31];
                Temp6_and_Next_ADDR_Data_29 <= {Temp6_and_Next_ADDR_Data_29[36:0], 1'b0};
                
                Slide_data_30 <= Temp6_and_Next_ADDR_Data_30[37:31];
                Temp6_and_Next_ADDR_Data_30 <= {Temp6_and_Next_ADDR_Data_30[36:0], 1'b0};
                
                Slide_data_31 <= Temp6_and_Next_ADDR_Data_31[37:31];
                Temp6_and_Next_ADDR_Data_31 <= {Temp6_and_Next_ADDR_Data_31[36:0], 1'b0};
                
                Slide_data_32 <= Temp6_and_Next_ADDR_Data_32[37:31];
                Temp6_and_Next_ADDR_Data_32 <= {Temp6_and_Next_ADDR_Data_32[36:0], 1'b0};
                
                Slide_data_33 <= Temp6_and_Next_ADDR_Data_33[37:31];
                Temp6_and_Next_ADDR_Data_33 <= {Temp6_and_Next_ADDR_Data_33[36:0], 1'b0};
                
                Slide_data_34 <= Temp6_and_Next_ADDR_Data_34[37:31];
                Temp6_and_Next_ADDR_Data_34 <= {Temp6_and_Next_ADDR_Data_34[36:0], 1'b0};
                
                Slide_data_35 <= Temp6_and_Next_ADDR_Data_35[37:31];
                Temp6_and_Next_ADDR_Data_35 <= {Temp6_and_Next_ADDR_Data_35[36:0], 1'b0};
                
                Slide_data_36 <= Temp6_and_Next_ADDR_Data_36[37:31];
                Temp6_and_Next_ADDR_Data_36 <= {Temp6_and_Next_ADDR_Data_36[36:0], 1'b0};
                
                Slide_data_37 <= Temp6_and_Next_ADDR_Data_37[37:31];
                Temp6_and_Next_ADDR_Data_37 <= {Temp6_and_Next_ADDR_Data_37[36:0], 1'b0};
                
                Slide_data_38 <= Temp6_and_Next_ADDR_Data_38[37:31];
                Temp6_and_Next_ADDR_Data_38 <= {Temp6_and_Next_ADDR_Data_38[36:0], 1'b0};
                
                Slide_data_39 <= Temp6_and_Next_ADDR_Data_39[37:31];
                Temp6_and_Next_ADDR_Data_39 <= {Temp6_and_Next_ADDR_Data_39[36:0], 1'b0};
                
                Slide_data_40 <= Temp6_and_Next_ADDR_Data_40[37:31];
                Temp6_and_Next_ADDR_Data_40 <= {Temp6_and_Next_ADDR_Data_40[36:0], 1'b0};
                
                Slide_data_41 <= Temp6_and_Next_ADDR_Data_41[37:31];
                Temp6_and_Next_ADDR_Data_41 <= {Temp6_and_Next_ADDR_Data_41[36:0], 1'b0};
                
                Slide_data_42 <= Temp6_and_Next_ADDR_Data_42[37:31];
                Temp6_and_Next_ADDR_Data_42 <= {Temp6_and_Next_ADDR_Data_42[36:0], 1'b0};
                
                Slide_data_43 <= Temp6_and_Next_ADDR_Data_43[37:31];
                Temp6_and_Next_ADDR_Data_43 <= {Temp6_and_Next_ADDR_Data_43[36:0], 1'b0};
                
                Slide_data_44 <= Temp6_and_Next_ADDR_Data_44[37:31];
                Temp6_and_Next_ADDR_Data_44 <= {Temp6_and_Next_ADDR_Data_44[36:0], 1'b0};
                
                Slide_data_45 <= Temp6_and_Next_ADDR_Data_45[37:31];
                Temp6_and_Next_ADDR_Data_45 <= {Temp6_and_Next_ADDR_Data_45[36:0], 1'b0};
                
                Slide_data_46 <= Temp6_and_Next_ADDR_Data_46[37:31];
                Temp6_and_Next_ADDR_Data_46 <= {Temp6_and_Next_ADDR_Data_46[36:0], 1'b0};
                
                Slide_data_47 <= Temp6_and_Next_ADDR_Data_47[37:31];
                Temp6_and_Next_ADDR_Data_47 <= {Temp6_and_Next_ADDR_Data_47[36:0], 1'b0};
                
                Slide_data_48 <= Temp6_and_Next_ADDR_Data_48[37:31];
                Temp6_and_Next_ADDR_Data_48 <= {Temp6_and_Next_ADDR_Data_48[36:0], 1'b0};
                
                Slide_data_49 <= Temp6_and_Next_ADDR_Data_49[37:31];
                Temp6_and_Next_ADDR_Data_49 <= {Temp6_and_Next_ADDR_Data_49[36:0], 1'b0};
                
                Slide_data_50 <= Temp6_and_Next_ADDR_Data_50[37:31];
                Temp6_and_Next_ADDR_Data_50 <= {Temp6_and_Next_ADDR_Data_50[36:0], 1'b0};
                
                Slide_data_51 <= Temp6_and_Next_ADDR_Data_51[37:31];
                Temp6_and_Next_ADDR_Data_51 <= {Temp6_and_Next_ADDR_Data_51[36:0], 1'b0};
                
                Slide_data_52 <= Temp6_and_Next_ADDR_Data_52[37:31];
                Temp6_and_Next_ADDR_Data_52 <= {Temp6_and_Next_ADDR_Data_52[36:0], 1'b0};
                
                Slide_data_53 <= Temp6_and_Next_ADDR_Data_53[37:31];
                Temp6_and_Next_ADDR_Data_53 <= {Temp6_and_Next_ADDR_Data_53[36:0], 1'b0};
                
                Slide_data_54 <= Temp6_and_Next_ADDR_Data_54[37:31];
                Temp6_and_Next_ADDR_Data_54 <= {Temp6_and_Next_ADDR_Data_54[36:0], 1'b0};
                
                Slide_data_55 <= Temp6_and_Next_ADDR_Data_55[37:31];
                Temp6_and_Next_ADDR_Data_55 <= {Temp6_and_Next_ADDR_Data_55[36:0], 1'b0};
                
                Slide_data_56 <= Temp6_and_Next_ADDR_Data_56[37:31];
                Temp6_and_Next_ADDR_Data_56 <= {Temp6_and_Next_ADDR_Data_56[36:0], 1'b0};
                
                Slide_data_57 <= Temp6_and_Next_ADDR_Data_57[37:31];
                Temp6_and_Next_ADDR_Data_57 <= {Temp6_and_Next_ADDR_Data_57[36:0], 1'b0};
                
                Slide_data_58 <= Temp6_and_Next_ADDR_Data_58[37:31];
                Temp6_and_Next_ADDR_Data_58 <= {Temp6_and_Next_ADDR_Data_58[36:0], 1'b0};
                
                Slide_data_59 <= Temp6_and_Next_ADDR_Data_59[37:31];
                Temp6_and_Next_ADDR_Data_59 <= {Temp6_and_Next_ADDR_Data_59[36:0], 1'b0};
                
                Slide_data_60 <= Temp6_and_Next_ADDR_Data_60[37:31];
                Temp6_and_Next_ADDR_Data_60 <= {Temp6_and_Next_ADDR_Data_60[36:0], 1'b0};
                
                Slide_data_61 <= Temp6_and_Next_ADDR_Data_61[37:31];
                Temp6_and_Next_ADDR_Data_61 <= {Temp6_and_Next_ADDR_Data_61[36:0], 1'b0};
                
                Slide_data_62 <= Temp6_and_Next_ADDR_Data_62[37:31];
                Temp6_and_Next_ADDR_Data_62 <= {Temp6_and_Next_ADDR_Data_62[36:0], 1'b0};
                
                Slide_data_63 <= Temp6_and_Next_ADDR_Data_63[37:31];
                Temp6_and_Next_ADDR_Data_63 <= {Temp6_and_Next_ADDR_Data_63[36:0], 1'b0};            
                if(cnt == 22)begin
                    Temp6_and_five_one_0 <= {Temp6_and_Next_ADDR_Data_0[36:31], padding_data[4:0]};
                    Temp6_and_five_one_1 <= {Temp6_and_Next_ADDR_Data_1[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_2 <= {Temp6_and_Next_ADDR_Data_2[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_3 <= {Temp6_and_Next_ADDR_Data_3[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_4 <= {Temp6_and_Next_ADDR_Data_4[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_5 <= {Temp6_and_Next_ADDR_Data_5[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_6 <= {Temp6_and_Next_ADDR_Data_6[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_7 <= {Temp6_and_Next_ADDR_Data_7[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_8 <= {Temp6_and_Next_ADDR_Data_8[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_9 <= {Temp6_and_Next_ADDR_Data_9[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_10 <= {Temp6_and_Next_ADDR_Data_10[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_11 <= {Temp6_and_Next_ADDR_Data_11[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_12 <= {Temp6_and_Next_ADDR_Data_12[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_13 <= {Temp6_and_Next_ADDR_Data_13[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_14 <= {Temp6_and_Next_ADDR_Data_14[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_15 <= {Temp6_and_Next_ADDR_Data_15[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_16 <= {Temp6_and_Next_ADDR_Data_16[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_17 <= {Temp6_and_Next_ADDR_Data_17[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_18 <= {Temp6_and_Next_ADDR_Data_18[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_19 <= {Temp6_and_Next_ADDR_Data_19[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_20 <= {Temp6_and_Next_ADDR_Data_20[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_21 <= {Temp6_and_Next_ADDR_Data_21[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_22 <= {Temp6_and_Next_ADDR_Data_22[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_23 <= {Temp6_and_Next_ADDR_Data_23[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_24 <= {Temp6_and_Next_ADDR_Data_24[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_25 <= {Temp6_and_Next_ADDR_Data_25[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_26 <= {Temp6_and_Next_ADDR_Data_26[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_27 <= {Temp6_and_Next_ADDR_Data_27[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_28 <= {Temp6_and_Next_ADDR_Data_28[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_29 <= {Temp6_and_Next_ADDR_Data_29[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_30 <= {Temp6_and_Next_ADDR_Data_30[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_31 <= {Temp6_and_Next_ADDR_Data_31[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_32 <= {Temp6_and_Next_ADDR_Data_32[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_33 <= {Temp6_and_Next_ADDR_Data_33[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_34 <= {Temp6_and_Next_ADDR_Data_34[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_35 <= {Temp6_and_Next_ADDR_Data_35[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_36 <= {Temp6_and_Next_ADDR_Data_36[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_37 <= {Temp6_and_Next_ADDR_Data_37[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_38 <= {Temp6_and_Next_ADDR_Data_38[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_39 <= {Temp6_and_Next_ADDR_Data_39[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_40 <= {Temp6_and_Next_ADDR_Data_40[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_41 <= {Temp6_and_Next_ADDR_Data_41[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_42 <= {Temp6_and_Next_ADDR_Data_42[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_43 <= {Temp6_and_Next_ADDR_Data_43[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_44 <= {Temp6_and_Next_ADDR_Data_44[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_45 <= {Temp6_and_Next_ADDR_Data_45[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_46 <= {Temp6_and_Next_ADDR_Data_46[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_47 <= {Temp6_and_Next_ADDR_Data_47[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_48 <= {Temp6_and_Next_ADDR_Data_48[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_49 <= {Temp6_and_Next_ADDR_Data_49[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_50 <= {Temp6_and_Next_ADDR_Data_50[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_51 <= {Temp6_and_Next_ADDR_Data_51[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_52 <= {Temp6_and_Next_ADDR_Data_52[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_53 <= {Temp6_and_Next_ADDR_Data_53[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_54 <= {Temp6_and_Next_ADDR_Data_54[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_55 <= {Temp6_and_Next_ADDR_Data_55[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_56 <= {Temp6_and_Next_ADDR_Data_56[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_57 <= {Temp6_and_Next_ADDR_Data_57[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_58 <= {Temp6_and_Next_ADDR_Data_58[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_59 <= {Temp6_and_Next_ADDR_Data_59[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_60 <= {Temp6_and_Next_ADDR_Data_60[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_61 <= {Temp6_and_Next_ADDR_Data_61[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_62 <= {Temp6_and_Next_ADDR_Data_62[36:31], padding_data[4:0]};        
                    Temp6_and_five_one_63 <= {Temp6_and_Next_ADDR_Data_63[36:31], padding_data[4:0]};        
                end
            end
            else if(cnt <= 27)begin
                Slide_data_0 <= Temp6_and_five_one_0[10:4];
                Temp6_and_five_one_0 <= {Temp6_and_five_one_0[9:0], 1'b0};
                
                Slide_data_1 <= Temp6_and_five_one_1[10:4];
                Temp6_and_five_one_1 <= {Temp6_and_five_one_1[9:0], 1'b0};       
                
                
                Slide_data_2 <= Temp6_and_five_one_2[10:4];
                Temp6_and_five_one_2 <= {Temp6_and_five_one_2[9:0], 1'b0};       
                
                
                Slide_data_3 <= Temp6_and_five_one_3[10:4];
                Temp6_and_five_one_3 <= {Temp6_and_five_one_3[9:0], 1'b0};       
                
                
                Slide_data_4 <= Temp6_and_five_one_4[10:4];
                Temp6_and_five_one_4 <= {Temp6_and_five_one_4[9:0], 1'b0};       
                
                
                Slide_data_5 <= Temp6_and_five_one_5[10:4];
                Temp6_and_five_one_5 <= {Temp6_and_five_one_5[9:0], 1'b0};       
                
                
                Slide_data_6 <= Temp6_and_five_one_6[10:4];
                Temp6_and_five_one_6 <= {Temp6_and_five_one_6[9:0], 1'b0};       
                
                
                Slide_data_7 <= Temp6_and_five_one_7[10:4];
                Temp6_and_five_one_7 <= {Temp6_and_five_one_7[9:0], 1'b0};       
                
                
                Slide_data_8 <= Temp6_and_five_one_8[10:4];
                Temp6_and_five_one_8 <= {Temp6_and_five_one_8[9:0], 1'b0};       
                
                
                Slide_data_9 <= Temp6_and_five_one_9[10:4];
                Temp6_and_five_one_9 <= {Temp6_and_five_one_9[9:0], 1'b0};       
                
                
                Slide_data_10 <= Temp6_and_five_one_10[10:4];
                Temp6_and_five_one_10 <= {Temp6_and_five_one_10[9:0], 1'b0};       
                
                
                Slide_data_11 <= Temp6_and_five_one_11[10:4];
                Temp6_and_five_one_11 <= {Temp6_and_five_one_11[9:0], 1'b0};       
                
                
                Slide_data_12 <= Temp6_and_five_one_12[10:4];
                Temp6_and_five_one_12 <= {Temp6_and_five_one_12[9:0], 1'b0};       
                
                
                Slide_data_13 <= Temp6_and_five_one_13[10:4];
                Temp6_and_five_one_13 <= {Temp6_and_five_one_13[9:0], 1'b0};       
                
                
                Slide_data_14 <= Temp6_and_five_one_14[10:4];
                Temp6_and_five_one_14 <= {Temp6_and_five_one_14[9:0], 1'b0};       
                
                
                Slide_data_15 <= Temp6_and_five_one_15[10:4];
                Temp6_and_five_one_15 <= {Temp6_and_five_one_15[9:0], 1'b0};       
                
                
                Slide_data_16 <= Temp6_and_five_one_16[10:4];
                Temp6_and_five_one_16 <= {Temp6_and_five_one_16[9:0], 1'b0};       
                
                
                Slide_data_17 <= Temp6_and_five_one_17[10:4];
                Temp6_and_five_one_17 <= {Temp6_and_five_one_17[9:0], 1'b0};       
                
                
                Slide_data_18 <= Temp6_and_five_one_18[10:4];
                Temp6_and_five_one_18 <= {Temp6_and_five_one_18[9:0], 1'b0};       
                
                
                Slide_data_19 <= Temp6_and_five_one_19[10:4];
                Temp6_and_five_one_19 <= {Temp6_and_five_one_19[9:0], 1'b0};       
                
                
                Slide_data_20 <= Temp6_and_five_one_20[10:4];
                Temp6_and_five_one_20 <= {Temp6_and_five_one_20[9:0], 1'b0};       
                
                
                Slide_data_21 <= Temp6_and_five_one_21[10:4];
                Temp6_and_five_one_21 <= {Temp6_and_five_one_21[9:0], 1'b0};       
                
                
                Slide_data_22 <= Temp6_and_five_one_22[10:4];
                Temp6_and_five_one_22 <= {Temp6_and_five_one_22[9:0], 1'b0};       
                
                
                Slide_data_23 <= Temp6_and_five_one_23[10:4];
                Temp6_and_five_one_23 <= {Temp6_and_five_one_23[9:0], 1'b0};       
                
                
                Slide_data_24 <= Temp6_and_five_one_24[10:4];
                Temp6_and_five_one_24 <= {Temp6_and_five_one_24[9:0], 1'b0};       
                
                
                Slide_data_25 <= Temp6_and_five_one_25[10:4];
                Temp6_and_five_one_25 <= {Temp6_and_five_one_25[9:0], 1'b0};       
                
                
                Slide_data_26 <= Temp6_and_five_one_26[10:4];
                Temp6_and_five_one_26 <= {Temp6_and_five_one_26[9:0], 1'b0};       
                
                
                Slide_data_27 <= Temp6_and_five_one_27[10:4];
                Temp6_and_five_one_27 <= {Temp6_and_five_one_27[9:0], 1'b0};       
                
                
                Slide_data_28 <= Temp6_and_five_one_28[10:4];
                Temp6_and_five_one_28 <= {Temp6_and_five_one_28[9:0], 1'b0};       
                
                
                Slide_data_29 <= Temp6_and_five_one_29[10:4];
                Temp6_and_five_one_29 <= {Temp6_and_five_one_29[9:0], 1'b0};       
                
                
                Slide_data_30 <= Temp6_and_five_one_30[10:4];
                Temp6_and_five_one_30 <= {Temp6_and_five_one_30[9:0], 1'b0};       
                
                
                Slide_data_31 <= Temp6_and_five_one_31[10:4];
                Temp6_and_five_one_31 <= {Temp6_and_five_one_31[9:0], 1'b0};       
                
                
                Slide_data_32 <= Temp6_and_five_one_32[10:4];
                Temp6_and_five_one_32 <= {Temp6_and_five_one_32[9:0], 1'b0};       
                
                
                Slide_data_33 <= Temp6_and_five_one_33[10:4];
                Temp6_and_five_one_33 <= {Temp6_and_five_one_33[9:0], 1'b0};       
                
                
                Slide_data_34 <= Temp6_and_five_one_34[10:4];
                Temp6_and_five_one_34 <= {Temp6_and_five_one_34[9:0], 1'b0};       
                
                
                Slide_data_35 <= Temp6_and_five_one_35[10:4];
                Temp6_and_five_one_35 <= {Temp6_and_five_one_35[9:0], 1'b0};       
                
                
                Slide_data_36 <= Temp6_and_five_one_36[10:4];
                Temp6_and_five_one_36 <= {Temp6_and_five_one_36[9:0], 1'b0};       
                
                
                Slide_data_37 <= Temp6_and_five_one_37[10:4];
                Temp6_and_five_one_37 <= {Temp6_and_five_one_37[9:0], 1'b0};       
                
                
                Slide_data_38 <= Temp6_and_five_one_38[10:4];
                Temp6_and_five_one_38 <= {Temp6_and_five_one_38[9:0], 1'b0};       
                
                
                Slide_data_39 <= Temp6_and_five_one_39[10:4];
                Temp6_and_five_one_39 <= {Temp6_and_five_one_39[9:0], 1'b0};       
                
                
                Slide_data_40 <= Temp6_and_five_one_40[10:4];
                Temp6_and_five_one_40 <= {Temp6_and_five_one_40[9:0], 1'b0};       
                
                
                Slide_data_41 <= Temp6_and_five_one_41[10:4];
                Temp6_and_five_one_41 <= {Temp6_and_five_one_41[9:0], 1'b0};       
                
                
                Slide_data_42 <= Temp6_and_five_one_42[10:4];
                Temp6_and_five_one_42 <= {Temp6_and_five_one_42[9:0], 1'b0};       
                
                
                Slide_data_43 <= Temp6_and_five_one_43[10:4];
                Temp6_and_five_one_43 <= {Temp6_and_five_one_43[9:0], 1'b0};       
                
                
                Slide_data_44 <= Temp6_and_five_one_44[10:4];
                Temp6_and_five_one_44 <= {Temp6_and_five_one_44[9:0], 1'b0};       
                
                
                Slide_data_45 <= Temp6_and_five_one_45[10:4];
                Temp6_and_five_one_45 <= {Temp6_and_five_one_45[9:0], 1'b0};       
                
                
                Slide_data_46 <= Temp6_and_five_one_46[10:4];
                Temp6_and_five_one_46 <= {Temp6_and_five_one_46[9:0], 1'b0};       
                
                
                Slide_data_47 <= Temp6_and_five_one_47[10:4];
                Temp6_and_five_one_47 <= {Temp6_and_five_one_47[9:0], 1'b0};       
                
                
                Slide_data_48 <= Temp6_and_five_one_48[10:4];
                Temp6_and_five_one_48 <= {Temp6_and_five_one_48[9:0], 1'b0};       
                
                
                Slide_data_49 <= Temp6_and_five_one_49[10:4];
                Temp6_and_five_one_49 <= {Temp6_and_five_one_49[9:0], 1'b0};       
                
                
                Slide_data_50 <= Temp6_and_five_one_50[10:4];
                Temp6_and_five_one_50 <= {Temp6_and_five_one_50[9:0], 1'b0};       
                
                
                Slide_data_51 <= Temp6_and_five_one_51[10:4];
                Temp6_and_five_one_51 <= {Temp6_and_five_one_51[9:0], 1'b0};       
                
                
                Slide_data_52 <= Temp6_and_five_one_52[10:4];
                Temp6_and_five_one_52 <= {Temp6_and_five_one_52[9:0], 1'b0};       
                
                
                Slide_data_53 <= Temp6_and_five_one_53[10:4];
                Temp6_and_five_one_53 <= {Temp6_and_five_one_53[9:0], 1'b0};       
                
                
                Slide_data_54 <= Temp6_and_five_one_54[10:4];
                Temp6_and_five_one_54 <= {Temp6_and_five_one_54[9:0], 1'b0};       
                
                
                Slide_data_55 <= Temp6_and_five_one_55[10:4];
                Temp6_and_five_one_55 <= {Temp6_and_five_one_55[9:0], 1'b0};       
                
                
                Slide_data_56 <= Temp6_and_five_one_56[10:4];
                Temp6_and_five_one_56 <= {Temp6_and_five_one_56[9:0], 1'b0};       
                
                
                Slide_data_57 <= Temp6_and_five_one_57[10:4];
                Temp6_and_five_one_57 <= {Temp6_and_five_one_57[9:0], 1'b0};       
                
                
                Slide_data_58 <= Temp6_and_five_one_58[10:4];
                Temp6_and_five_one_58 <= {Temp6_and_five_one_58[9:0], 1'b0};       
                
                
                Slide_data_59 <= Temp6_and_five_one_59[10:4];
                Temp6_and_five_one_59 <= {Temp6_and_five_one_59[9:0], 1'b0};       
                
                
                Slide_data_60 <= Temp6_and_five_one_60[10:4];
                Temp6_and_five_one_60 <= {Temp6_and_five_one_60[9:0], 1'b0};       
                
                
                Slide_data_61 <= Temp6_and_five_one_61[10:4];
                Temp6_and_five_one_61 <= {Temp6_and_five_one_61[9:0], 1'b0};       
                
                
                Slide_data_62 <= Temp6_and_five_one_62[10:4];
                Temp6_and_five_one_62 <= {Temp6_and_five_one_62[9:0], 1'b0};       
                
                
                Slide_data_63 <= Temp6_and_five_one_63[10:4];
                Temp6_and_five_one_63 <= {Temp6_and_five_one_63[9:0], 1'b0};       
            end
          else begin
            padding_data <= 0;
            
            Slide_data_0 <= 0;
            Temp6_0      <= 0;
            Pad_and_ADDR1_Temp_0 <= 0;
            Temp6_and_Next_ADDR_Data_0 <= 0;
            Temp6_and_five_one_0 <= 0;
            
            Slide_data_1 <= 0;
                Temp6_1      <= 0;
                Pad_and_ADDR1_Temp_1 <= 0;
                Temp6_and_Next_ADDR_Data_1 <= 0;
                Temp6_and_five_one_1 <= 0;       
                
                
                Slide_data_2 <= 0;
                Temp6_2      <= 0;
                Pad_and_ADDR1_Temp_2 <= 0;
                Temp6_and_Next_ADDR_Data_2 <= 0;
                Temp6_and_five_one_2 <= 0;       
                
                
                Slide_data_3 <= 0;
                Temp6_3      <= 0;
                Pad_and_ADDR1_Temp_3 <= 0;
                Temp6_and_Next_ADDR_Data_3 <= 0;
                Temp6_and_five_one_3 <= 0;       
                
                
                Slide_data_4 <= 0;
                Temp6_4      <= 0;
                Pad_and_ADDR1_Temp_4 <= 0;
                Temp6_and_Next_ADDR_Data_4 <= 0;
                Temp6_and_five_one_4 <= 0;       
                
                
                Slide_data_5 <= 0;
                Temp6_5      <= 0;
                Pad_and_ADDR1_Temp_5 <= 0;
                Temp6_and_Next_ADDR_Data_5 <= 0;
                Temp6_and_five_one_5 <= 0;       
                
                
                Slide_data_6 <= 0;
                Temp6_6      <= 0;
                Pad_and_ADDR1_Temp_6 <= 0;
                Temp6_and_Next_ADDR_Data_6 <= 0;
                Temp6_and_five_one_6 <= 0;       
                
                
                Slide_data_7 <= 0;
                Temp6_7      <= 0;
                Pad_and_ADDR1_Temp_7 <= 0;
                Temp6_and_Next_ADDR_Data_7 <= 0;
                Temp6_and_five_one_7 <= 0;       
                
                
                Slide_data_8 <= 0;
                Temp6_8      <= 0;
                Pad_and_ADDR1_Temp_8 <= 0;
                Temp6_and_Next_ADDR_Data_8 <= 0;
                Temp6_and_five_one_8 <= 0;       
                
                
                Slide_data_9 <= 0;
                Temp6_9      <= 0;
                Pad_and_ADDR1_Temp_9 <= 0;
                Temp6_and_Next_ADDR_Data_9 <= 0;
                Temp6_and_five_one_9 <= 0;       
                
                
                Slide_data_10 <= 0;
                Temp6_10      <= 0;
                Pad_and_ADDR1_Temp_10 <= 0;
                Temp6_and_Next_ADDR_Data_10 <= 0;
                Temp6_and_five_one_10 <= 0;       
                
                
                Slide_data_11 <= 0;
                Temp6_11      <= 0;
                Pad_and_ADDR1_Temp_11 <= 0;
                Temp6_and_Next_ADDR_Data_11 <= 0;
                Temp6_and_five_one_11 <= 0;       
                
                
                Slide_data_12 <= 0;
                Temp6_12      <= 0;
                Pad_and_ADDR1_Temp_12 <= 0;
                Temp6_and_Next_ADDR_Data_12 <= 0;
                Temp6_and_five_one_12 <= 0;       
                
                
                Slide_data_13 <= 0;
                Temp6_13      <= 0;
                Pad_and_ADDR1_Temp_13 <= 0;
                Temp6_and_Next_ADDR_Data_13 <= 0;
                Temp6_and_five_one_13 <= 0;       
                
                
                Slide_data_14 <= 0;
                Temp6_14      <= 0;
                Pad_and_ADDR1_Temp_14 <= 0;
                Temp6_and_Next_ADDR_Data_14 <= 0;
                Temp6_and_five_one_14 <= 0;       
                
                
                Slide_data_15 <= 0;
                Temp6_15      <= 0;
                Pad_and_ADDR1_Temp_15 <= 0;
                Temp6_and_Next_ADDR_Data_15 <= 0;
                Temp6_and_five_one_15 <= 0;       
                
                
                Slide_data_16 <= 0;
                Temp6_16      <= 0;
                Pad_and_ADDR1_Temp_16 <= 0;
                Temp6_and_Next_ADDR_Data_16 <= 0;
                Temp6_and_five_one_16 <= 0;       
                
                
                Slide_data_17 <= 0;
                Temp6_17      <= 0;
                Pad_and_ADDR1_Temp_17 <= 0;
                Temp6_and_Next_ADDR_Data_17 <= 0;
                Temp6_and_five_one_17 <= 0;       
                
                
                Slide_data_18 <= 0;
                Temp6_18      <= 0;
                Pad_and_ADDR1_Temp_18 <= 0;
                Temp6_and_Next_ADDR_Data_18 <= 0;
                Temp6_and_five_one_18 <= 0;       
                
                
                Slide_data_19 <= 0;
                Temp6_19      <= 0;
                Pad_and_ADDR1_Temp_19 <= 0;
                Temp6_and_Next_ADDR_Data_19 <= 0;
                Temp6_and_five_one_19 <= 0;       
                
                
                Slide_data_20 <= 0;
                Temp6_20      <= 0;
                Pad_and_ADDR1_Temp_20 <= 0;
                Temp6_and_Next_ADDR_Data_20 <= 0;
                Temp6_and_five_one_20 <= 0;       
                
                
                Slide_data_21 <= 0;
                Temp6_21      <= 0;
                Pad_and_ADDR1_Temp_21 <= 0;
                Temp6_and_Next_ADDR_Data_21 <= 0;
                Temp6_and_five_one_21 <= 0;       
                
                
                Slide_data_22 <= 0;
                Temp6_22      <= 0;
                Pad_and_ADDR1_Temp_22 <= 0;
                Temp6_and_Next_ADDR_Data_22 <= 0;
                Temp6_and_five_one_22 <= 0;       
                
                
                Slide_data_23 <= 0;
                Temp6_23      <= 0;
                Pad_and_ADDR1_Temp_23 <= 0;
                Temp6_and_Next_ADDR_Data_23 <= 0;
                Temp6_and_five_one_23 <= 0;       
                
                
                Slide_data_24 <= 0;
                Temp6_24      <= 0;
                Pad_and_ADDR1_Temp_24 <= 0;
                Temp6_and_Next_ADDR_Data_24 <= 0;
                Temp6_and_five_one_24 <= 0;       
                
                
                Slide_data_25 <= 0;
                Temp6_25      <= 0;
                Pad_and_ADDR1_Temp_25 <= 0;
                Temp6_and_Next_ADDR_Data_25 <= 0;
                Temp6_and_five_one_25 <= 0;       
                
                
                Slide_data_26 <= 0;
                Temp6_26      <= 0;
                Pad_and_ADDR1_Temp_26 <= 0;
                Temp6_and_Next_ADDR_Data_26 <= 0;
                Temp6_and_five_one_26 <= 0;       
                
                
                Slide_data_27 <= 0;
                Temp6_27      <= 0;
                Pad_and_ADDR1_Temp_27 <= 0;
                Temp6_and_Next_ADDR_Data_27 <= 0;
                Temp6_and_five_one_27 <= 0;       
                
                
                Slide_data_28 <= 0;
                Temp6_28      <= 0;
                Pad_and_ADDR1_Temp_28 <= 0;
                Temp6_and_Next_ADDR_Data_28 <= 0;
                Temp6_and_five_one_28 <= 0;       
                
                
                Slide_data_29 <= 0;
                Temp6_29      <= 0;
                Pad_and_ADDR1_Temp_29 <= 0;
                Temp6_and_Next_ADDR_Data_29 <= 0;
                Temp6_and_five_one_29 <= 0;       
                
                
                Slide_data_30 <= 0;
                Temp6_30      <= 0;
                Pad_and_ADDR1_Temp_30 <= 0;
                Temp6_and_Next_ADDR_Data_30 <= 0;
                Temp6_and_five_one_30 <= 0;       
                
                
                Slide_data_31 <= 0;
                Temp6_31      <= 0;
                Pad_and_ADDR1_Temp_31 <= 0;
                Temp6_and_Next_ADDR_Data_31 <= 0;
                Temp6_and_five_one_31 <= 0;       
                
                
                Slide_data_32 <= 0;
                Temp6_32      <= 0;
                Pad_and_ADDR1_Temp_32 <= 0;
                Temp6_and_Next_ADDR_Data_32 <= 0;
                Temp6_and_five_one_32 <= 0;       
                
                
                Slide_data_33 <= 0;
                Temp6_33      <= 0;
                Pad_and_ADDR1_Temp_33 <= 0;
                Temp6_and_Next_ADDR_Data_33 <= 0;
                Temp6_and_five_one_33 <= 0;       
                
                
                Slide_data_34 <= 0;
                Temp6_34      <= 0;
                Pad_and_ADDR1_Temp_34 <= 0;
                Temp6_and_Next_ADDR_Data_34 <= 0;
                Temp6_and_five_one_34 <= 0;       
                
                
                Slide_data_35 <= 0;
                Temp6_35      <= 0;
                Pad_and_ADDR1_Temp_35 <= 0;
                Temp6_and_Next_ADDR_Data_35 <= 0;
                Temp6_and_five_one_35 <= 0;       
                
                
                Slide_data_36 <= 0;
                Temp6_36      <= 0;
                Pad_and_ADDR1_Temp_36 <= 0;
                Temp6_and_Next_ADDR_Data_36 <= 0;
                Temp6_and_five_one_36 <= 0;       
                
                
                Slide_data_37 <= 0;
                Temp6_37      <= 0;
                Pad_and_ADDR1_Temp_37 <= 0;
                Temp6_and_Next_ADDR_Data_37 <= 0;
                Temp6_and_five_one_37 <= 0;       
                
                
                Slide_data_38 <= 0;
                Temp6_38      <= 0;
                Pad_and_ADDR1_Temp_38 <= 0;
                Temp6_and_Next_ADDR_Data_38 <= 0;
                Temp6_and_five_one_38 <= 0;       
                
                
                Slide_data_39 <= 0;
                Temp6_39      <= 0;
                Pad_and_ADDR1_Temp_39 <= 0;
                Temp6_and_Next_ADDR_Data_39 <= 0;
                Temp6_and_five_one_39 <= 0;       
                
                
                Slide_data_40 <= 0;
                Temp6_40      <= 0;
                Pad_and_ADDR1_Temp_40 <= 0;
                Temp6_and_Next_ADDR_Data_40 <= 0;
                Temp6_and_five_one_40 <= 0;       
                
                
                Slide_data_41 <= 0;
                Temp6_41      <= 0;
                Pad_and_ADDR1_Temp_41 <= 0;
                Temp6_and_Next_ADDR_Data_41 <= 0;
                Temp6_and_five_one_41 <= 0;       
                
                
                Slide_data_42 <= 0;
                Temp6_42      <= 0;
                Pad_and_ADDR1_Temp_42 <= 0;
                Temp6_and_Next_ADDR_Data_42 <= 0;
                Temp6_and_five_one_42 <= 0;       
                
                
                Slide_data_43 <= 0;
                Temp6_43      <= 0;
                Pad_and_ADDR1_Temp_43 <= 0;
                Temp6_and_Next_ADDR_Data_43 <= 0;
                Temp6_and_five_one_43 <= 0;       
                
                
                Slide_data_44 <= 0;
                Temp6_44      <= 0;
                Pad_and_ADDR1_Temp_44 <= 0;
                Temp6_and_Next_ADDR_Data_44 <= 0;
                Temp6_and_five_one_44 <= 0;       
                
                
                Slide_data_45 <= 0;
                Temp6_45      <= 0;
                Pad_and_ADDR1_Temp_45 <= 0;
                Temp6_and_Next_ADDR_Data_45 <= 0;
                Temp6_and_five_one_45 <= 0;       
                
                
                Slide_data_46 <= 0;
                Temp6_46      <= 0;
                Pad_and_ADDR1_Temp_46 <= 0;
                Temp6_and_Next_ADDR_Data_46 <= 0;
                Temp6_and_five_one_46 <= 0;       
                
                
                Slide_data_47 <= 0;
                Temp6_47      <= 0;
                Pad_and_ADDR1_Temp_47 <= 0;
                Temp6_and_Next_ADDR_Data_47 <= 0;
                Temp6_and_five_one_47 <= 0;       
                
                
                Slide_data_48 <= 0;
                Temp6_48      <= 0;
                Pad_and_ADDR1_Temp_48 <= 0;
                Temp6_and_Next_ADDR_Data_48 <= 0;
                Temp6_and_five_one_48 <= 0;       
                
                
                Slide_data_49 <= 0;
                Temp6_49      <= 0;
                Pad_and_ADDR1_Temp_49 <= 0;
                Temp6_and_Next_ADDR_Data_49 <= 0;
                Temp6_and_five_one_49 <= 0;       
                
                
                Slide_data_50 <= 0;
                Temp6_50      <= 0;
                Pad_and_ADDR1_Temp_50 <= 0;
                Temp6_and_Next_ADDR_Data_50 <= 0;
                Temp6_and_five_one_50 <= 0;       
                
                
                Slide_data_51 <= 0;
                Temp6_51      <= 0;
                Pad_and_ADDR1_Temp_51 <= 0;
                Temp6_and_Next_ADDR_Data_51 <= 0;
                Temp6_and_five_one_51 <= 0;       
                
                
                Slide_data_52 <= 0;
                Temp6_52      <= 0;
                Pad_and_ADDR1_Temp_52 <= 0;
                Temp6_and_Next_ADDR_Data_52 <= 0;
                Temp6_and_five_one_52 <= 0;       
                
                
                Slide_data_53 <= 0;
                Temp6_53      <= 0;
                Pad_and_ADDR1_Temp_53 <= 0;
                Temp6_and_Next_ADDR_Data_53 <= 0;
                Temp6_and_five_one_53 <= 0;       
                
                
                Slide_data_54 <= 0;
                Temp6_54      <= 0;
                Pad_and_ADDR1_Temp_54 <= 0;
                Temp6_and_Next_ADDR_Data_54 <= 0;
                Temp6_and_five_one_54 <= 0;       
                
                
                Slide_data_55 <= 0;
                Temp6_55      <= 0;
                Pad_and_ADDR1_Temp_55 <= 0;
                Temp6_and_Next_ADDR_Data_55 <= 0;
                Temp6_and_five_one_55 <= 0;       
                
                
                Slide_data_56 <= 0;
                Temp6_56      <= 0;
                Pad_and_ADDR1_Temp_56 <= 0;
                Temp6_and_Next_ADDR_Data_56 <= 0;
                Temp6_and_five_one_56 <= 0;       
                
                
                Slide_data_57 <= 0;
                Temp6_57      <= 0;
                Pad_and_ADDR1_Temp_57 <= 0;
                Temp6_and_Next_ADDR_Data_57 <= 0;
                Temp6_and_five_one_57 <= 0;       
                
                
                Slide_data_58 <= 0;
                Temp6_58      <= 0;
                Pad_and_ADDR1_Temp_58 <= 0;
                Temp6_and_Next_ADDR_Data_58 <= 0;
                Temp6_and_five_one_58 <= 0;       
                
                
                Slide_data_59 <= 0;
                Temp6_59      <= 0;
                Pad_and_ADDR1_Temp_59 <= 0;
                Temp6_and_Next_ADDR_Data_59 <= 0;
                Temp6_and_five_one_59 <= 0;       
                
                
                Slide_data_60 <= 0;
                Temp6_60      <= 0;
                Pad_and_ADDR1_Temp_60 <= 0;
                Temp6_and_Next_ADDR_Data_60 <= 0;
                Temp6_and_five_one_60 <= 0;       
                
                
                Slide_data_61 <= 0;
                Temp6_61      <= 0;
                Pad_and_ADDR1_Temp_61 <= 0;
                Temp6_and_Next_ADDR_Data_61 <= 0;
                Temp6_and_five_one_61 <= 0;       
                
                
                Slide_data_62 <= 0;
                Temp6_62      <= 0;
                Pad_and_ADDR1_Temp_62 <= 0;
                Temp6_and_Next_ADDR_Data_62 <= 0;
                Temp6_and_five_one_62 <= 0;       
                
                
                Slide_data_63 <= 0;
                Temp6_63      <= 0;
                Pad_and_ADDR1_Temp_63 <= 0;
                Temp6_and_Next_ADDR_Data_63 <= 0;
                Temp6_and_five_one_63 <= 0;              
          end
        end
     end
end





endmodule
