`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/05/08 09:38:37
// Design Name: 
// Module Name: PE_Array_B5
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module PE_Array_B5(
    input                       clk,
    input                       rst_n,
    input               [63:0]  new_weight_val,
    input               [6:0]   w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7, w_8, w_9, w_10, w_11, w_12, w_13, w_14, w_15,
                                w_16, w_17, w_18, w_19, w_20, w_21, w_22, w_23, w_24, w_25, w_26, w_27, w_28, w_29, w_30, w_31,
    input   wire        [6:0]   Slide_data_0, Slide_data_1, Slide_data_2, Slide_data_3, Slide_data_4, Slide_data_5, Slide_data_6, Slide_data_7,
                                Slide_data_8, Slide_data_9, Slide_data_10, Slide_data_11, Slide_data_12, Slide_data_13, Slide_data_14, Slide_data_15,
                                Slide_data_16, Slide_data_17, Slide_data_18, Slide_data_19, Slide_data_20, Slide_data_21, Slide_data_22, Slide_data_23, 
                                Slide_data_24, Slide_data_25, Slide_data_26, Slide_data_27, Slide_data_28, Slide_data_29, Slide_data_30, Slide_data_31,
    output  wire signed [8:0]   o_0, o_1, o_2, o_3, o_4, o_5, o_6, o_7, o_8, o_9, o_10, o_11, o_12, o_13, o_14, o_15,
                                o_16, o_17, o_18, o_19, o_20, o_21, o_22, o_23, o_24, o_25, o_26, o_27, o_28, o_29, o_30, o_31, 
                                o_32, o_33, o_34, o_35, o_36, o_37, o_38, o_39, o_40, o_41, o_42, o_43, o_44, o_45, o_46, o_47, 
                                o_48, o_49, o_50, o_51, o_52, o_53, o_54, o_55, o_56, o_57, o_58, o_59, o_60, o_61, o_62, o_63,
    output  wire                o_0_val  
);

wire    [6:0]           in_data_to_next_pe_0_0, in_data_to_next_pe_0_1, in_data_to_next_pe_0_2, in_data_to_next_pe_0_3,  
                        in_data_to_next_pe_0_4, in_data_to_next_pe_0_5, in_data_to_next_pe_0_6, in_data_to_next_pe_0_7,
                        in_data_to_next_pe_0_8, in_data_to_next_pe_0_9, in_data_to_next_pe_0_10, in_data_to_next_pe_0_11,
                        in_data_to_next_pe_0_12, in_data_to_next_pe_0_13, in_data_to_next_pe_0_14, in_data_to_next_pe_0_15,
                        in_data_to_next_pe_0_16, in_data_to_next_pe_0_17, in_data_to_next_pe_0_18, in_data_to_next_pe_0_19, 
                        in_data_to_next_pe_0_20, in_data_to_next_pe_0_21, in_data_to_next_pe_0_22, in_data_to_next_pe_0_23, 
                        in_data_to_next_pe_0_24, in_data_to_next_pe_0_25, in_data_to_next_pe_0_26, in_data_to_next_pe_0_27, 
                        in_data_to_next_pe_0_28, in_data_to_next_pe_0_29, in_data_to_next_pe_0_30, in_data_to_next_pe_0_31,
                        
                        in_data_to_next_pe_1_0, in_data_to_next_pe_1_1, in_data_to_next_pe_1_2, in_data_to_next_pe_1_3,  
                        in_data_to_next_pe_1_4, in_data_to_next_pe_1_5, in_data_to_next_pe_1_6, in_data_to_next_pe_1_7,
                        in_data_to_next_pe_1_8, in_data_to_next_pe_1_9, in_data_to_next_pe_1_10, in_data_to_next_pe_1_11,
                        in_data_to_next_pe_1_12, in_data_to_next_pe_1_13, in_data_to_next_pe_1_14, in_data_to_next_pe_1_15,
                        in_data_to_next_pe_1_16, in_data_to_next_pe_1_17, in_data_to_next_pe_1_18, in_data_to_next_pe_1_19, 
                        in_data_to_next_pe_1_20, in_data_to_next_pe_1_21, in_data_to_next_pe_1_22, in_data_to_next_pe_1_23, 
                        in_data_to_next_pe_1_24, in_data_to_next_pe_1_25, in_data_to_next_pe_1_26, in_data_to_next_pe_1_27, 
                        in_data_to_next_pe_1_28, in_data_to_next_pe_1_29, in_data_to_next_pe_1_30, in_data_to_next_pe_1_31, 
                        
                        
                        in_data_to_next_pe_2_0, in_data_to_next_pe_2_1, in_data_to_next_pe_2_2, in_data_to_next_pe_2_3,  
                        in_data_to_next_pe_2_4, in_data_to_next_pe_2_5, in_data_to_next_pe_2_6, in_data_to_next_pe_2_7,
                        in_data_to_next_pe_2_8, in_data_to_next_pe_2_9, in_data_to_next_pe_2_10, in_data_to_next_pe_2_11,
                        in_data_to_next_pe_2_12, in_data_to_next_pe_2_13, in_data_to_next_pe_2_14, in_data_to_next_pe_2_15,
                        in_data_to_next_pe_2_16, in_data_to_next_pe_2_17, in_data_to_next_pe_2_18, in_data_to_next_pe_2_19, 
                        in_data_to_next_pe_2_20, in_data_to_next_pe_2_21, in_data_to_next_pe_2_22, in_data_to_next_pe_2_23, 
                        in_data_to_next_pe_2_24, in_data_to_next_pe_2_25, in_data_to_next_pe_2_26, in_data_to_next_pe_2_27, 
                        in_data_to_next_pe_2_28, in_data_to_next_pe_2_29, in_data_to_next_pe_2_30, in_data_to_next_pe_2_31, 
                        
                        
                        in_data_to_next_pe_3_0, in_data_to_next_pe_3_1, in_data_to_next_pe_3_2, in_data_to_next_pe_3_3,  
                        in_data_to_next_pe_3_4, in_data_to_next_pe_3_5, in_data_to_next_pe_3_6, in_data_to_next_pe_3_7,
                        in_data_to_next_pe_3_8, in_data_to_next_pe_3_9, in_data_to_next_pe_3_10, in_data_to_next_pe_3_11,
                        in_data_to_next_pe_3_12, in_data_to_next_pe_3_13, in_data_to_next_pe_3_14, in_data_to_next_pe_3_15,
                        in_data_to_next_pe_3_16, in_data_to_next_pe_3_17, in_data_to_next_pe_3_18, in_data_to_next_pe_3_19, 
                        in_data_to_next_pe_3_20, in_data_to_next_pe_3_21, in_data_to_next_pe_3_22, in_data_to_next_pe_3_23, 
                        in_data_to_next_pe_3_24, in_data_to_next_pe_3_25, in_data_to_next_pe_3_26, in_data_to_next_pe_3_27, 
                        in_data_to_next_pe_3_28, in_data_to_next_pe_3_29, in_data_to_next_pe_3_30, in_data_to_next_pe_3_31, 
                        
                        
                        in_data_to_next_pe_4_0, in_data_to_next_pe_4_1, in_data_to_next_pe_4_2, in_data_to_next_pe_4_3,  
                        in_data_to_next_pe_4_4, in_data_to_next_pe_4_5, in_data_to_next_pe_4_6, in_data_to_next_pe_4_7,
                        in_data_to_next_pe_4_8, in_data_to_next_pe_4_9, in_data_to_next_pe_4_10, in_data_to_next_pe_4_11,
                        in_data_to_next_pe_4_12, in_data_to_next_pe_4_13, in_data_to_next_pe_4_14, in_data_to_next_pe_4_15,
                        in_data_to_next_pe_4_16, in_data_to_next_pe_4_17, in_data_to_next_pe_4_18, in_data_to_next_pe_4_19, 
                        in_data_to_next_pe_4_20, in_data_to_next_pe_4_21, in_data_to_next_pe_4_22, in_data_to_next_pe_4_23, 
                        in_data_to_next_pe_4_24, in_data_to_next_pe_4_25, in_data_to_next_pe_4_26, in_data_to_next_pe_4_27, 
                        in_data_to_next_pe_4_28, in_data_to_next_pe_4_29, in_data_to_next_pe_4_30, in_data_to_next_pe_4_31, 
                        
                        
                        in_data_to_next_pe_5_0, in_data_to_next_pe_5_1, in_data_to_next_pe_5_2, in_data_to_next_pe_5_3,  
                        in_data_to_next_pe_5_4, in_data_to_next_pe_5_5, in_data_to_next_pe_5_6, in_data_to_next_pe_5_7,
                        in_data_to_next_pe_5_8, in_data_to_next_pe_5_9, in_data_to_next_pe_5_10, in_data_to_next_pe_5_11,
                        in_data_to_next_pe_5_12, in_data_to_next_pe_5_13, in_data_to_next_pe_5_14, in_data_to_next_pe_5_15,
                        in_data_to_next_pe_5_16, in_data_to_next_pe_5_17, in_data_to_next_pe_5_18, in_data_to_next_pe_5_19, 
                        in_data_to_next_pe_5_20, in_data_to_next_pe_5_21, in_data_to_next_pe_5_22, in_data_to_next_pe_5_23, 
                        in_data_to_next_pe_5_24, in_data_to_next_pe_5_25, in_data_to_next_pe_5_26, in_data_to_next_pe_5_27, 
                        in_data_to_next_pe_5_28, in_data_to_next_pe_5_29, in_data_to_next_pe_5_30, in_data_to_next_pe_5_31, 
                        
                        
                        in_data_to_next_pe_6_0, in_data_to_next_pe_6_1, in_data_to_next_pe_6_2, in_data_to_next_pe_6_3,  
                        in_data_to_next_pe_6_4, in_data_to_next_pe_6_5, in_data_to_next_pe_6_6, in_data_to_next_pe_6_7,
                        in_data_to_next_pe_6_8, in_data_to_next_pe_6_9, in_data_to_next_pe_6_10, in_data_to_next_pe_6_11,
                        in_data_to_next_pe_6_12, in_data_to_next_pe_6_13, in_data_to_next_pe_6_14, in_data_to_next_pe_6_15,
                        in_data_to_next_pe_6_16, in_data_to_next_pe_6_17, in_data_to_next_pe_6_18, in_data_to_next_pe_6_19, 
                        in_data_to_next_pe_6_20, in_data_to_next_pe_6_21, in_data_to_next_pe_6_22, in_data_to_next_pe_6_23, 
                        in_data_to_next_pe_6_24, in_data_to_next_pe_6_25, in_data_to_next_pe_6_26, in_data_to_next_pe_6_27, 
                        in_data_to_next_pe_6_28, in_data_to_next_pe_6_29, in_data_to_next_pe_6_30, in_data_to_next_pe_6_31, 
                        
                        
                        in_data_to_next_pe_7_0, in_data_to_next_pe_7_1, in_data_to_next_pe_7_2, in_data_to_next_pe_7_3,  
                        in_data_to_next_pe_7_4, in_data_to_next_pe_7_5, in_data_to_next_pe_7_6, in_data_to_next_pe_7_7,
                        in_data_to_next_pe_7_8, in_data_to_next_pe_7_9, in_data_to_next_pe_7_10, in_data_to_next_pe_7_11,
                        in_data_to_next_pe_7_12, in_data_to_next_pe_7_13, in_data_to_next_pe_7_14, in_data_to_next_pe_7_15,
                        in_data_to_next_pe_7_16, in_data_to_next_pe_7_17, in_data_to_next_pe_7_18, in_data_to_next_pe_7_19, 
                        in_data_to_next_pe_7_20, in_data_to_next_pe_7_21, in_data_to_next_pe_7_22, in_data_to_next_pe_7_23, 
                        in_data_to_next_pe_7_24, in_data_to_next_pe_7_25, in_data_to_next_pe_7_26, in_data_to_next_pe_7_27, 
                        in_data_to_next_pe_7_28, in_data_to_next_pe_7_29, in_data_to_next_pe_7_30, in_data_to_next_pe_7_31, 
                        
                        
                        in_data_to_next_pe_8_0, in_data_to_next_pe_8_1, in_data_to_next_pe_8_2, in_data_to_next_pe_8_3,  
                        in_data_to_next_pe_8_4, in_data_to_next_pe_8_5, in_data_to_next_pe_8_6, in_data_to_next_pe_8_7,
                        in_data_to_next_pe_8_8, in_data_to_next_pe_8_9, in_data_to_next_pe_8_10, in_data_to_next_pe_8_11,
                        in_data_to_next_pe_8_12, in_data_to_next_pe_8_13, in_data_to_next_pe_8_14, in_data_to_next_pe_8_15,
                        in_data_to_next_pe_8_16, in_data_to_next_pe_8_17, in_data_to_next_pe_8_18, in_data_to_next_pe_8_19, 
                        in_data_to_next_pe_8_20, in_data_to_next_pe_8_21, in_data_to_next_pe_8_22, in_data_to_next_pe_8_23, 
                        in_data_to_next_pe_8_24, in_data_to_next_pe_8_25, in_data_to_next_pe_8_26, in_data_to_next_pe_8_27, 
                        in_data_to_next_pe_8_28, in_data_to_next_pe_8_29, in_data_to_next_pe_8_30, in_data_to_next_pe_8_31, 
                        
                        
                        in_data_to_next_pe_9_0, in_data_to_next_pe_9_1, in_data_to_next_pe_9_2, in_data_to_next_pe_9_3,  
                        in_data_to_next_pe_9_4, in_data_to_next_pe_9_5, in_data_to_next_pe_9_6, in_data_to_next_pe_9_7,
                        in_data_to_next_pe_9_8, in_data_to_next_pe_9_9, in_data_to_next_pe_9_10, in_data_to_next_pe_9_11,
                        in_data_to_next_pe_9_12, in_data_to_next_pe_9_13, in_data_to_next_pe_9_14, in_data_to_next_pe_9_15,
                        in_data_to_next_pe_9_16, in_data_to_next_pe_9_17, in_data_to_next_pe_9_18, in_data_to_next_pe_9_19, 
                        in_data_to_next_pe_9_20, in_data_to_next_pe_9_21, in_data_to_next_pe_9_22, in_data_to_next_pe_9_23, 
                        in_data_to_next_pe_9_24, in_data_to_next_pe_9_25, in_data_to_next_pe_9_26, in_data_to_next_pe_9_27, 
                        in_data_to_next_pe_9_28, in_data_to_next_pe_9_29, in_data_to_next_pe_9_30, in_data_to_next_pe_9_31, 
                        
                        
                        in_data_to_next_pe_10_0, in_data_to_next_pe_10_1, in_data_to_next_pe_10_2, in_data_to_next_pe_10_3,  
                        in_data_to_next_pe_10_4, in_data_to_next_pe_10_5, in_data_to_next_pe_10_6, in_data_to_next_pe_10_7,
                        in_data_to_next_pe_10_8, in_data_to_next_pe_10_9, in_data_to_next_pe_10_10, in_data_to_next_pe_10_11,
                        in_data_to_next_pe_10_12, in_data_to_next_pe_10_13, in_data_to_next_pe_10_14, in_data_to_next_pe_10_15,
                        in_data_to_next_pe_10_16, in_data_to_next_pe_10_17, in_data_to_next_pe_10_18, in_data_to_next_pe_10_19, 
                        in_data_to_next_pe_10_20, in_data_to_next_pe_10_21, in_data_to_next_pe_10_22, in_data_to_next_pe_10_23, 
                        in_data_to_next_pe_10_24, in_data_to_next_pe_10_25, in_data_to_next_pe_10_26, in_data_to_next_pe_10_27, 
                        in_data_to_next_pe_10_28, in_data_to_next_pe_10_29, in_data_to_next_pe_10_30, in_data_to_next_pe_10_31, 
                        
                        
                        in_data_to_next_pe_11_0, in_data_to_next_pe_11_1, in_data_to_next_pe_11_2, in_data_to_next_pe_11_3,  
                        in_data_to_next_pe_11_4, in_data_to_next_pe_11_5, in_data_to_next_pe_11_6, in_data_to_next_pe_11_7,
                        in_data_to_next_pe_11_8, in_data_to_next_pe_11_9, in_data_to_next_pe_11_10, in_data_to_next_pe_11_11,
                        in_data_to_next_pe_11_12, in_data_to_next_pe_11_13, in_data_to_next_pe_11_14, in_data_to_next_pe_11_15,
                        in_data_to_next_pe_11_16, in_data_to_next_pe_11_17, in_data_to_next_pe_11_18, in_data_to_next_pe_11_19, 
                        in_data_to_next_pe_11_20, in_data_to_next_pe_11_21, in_data_to_next_pe_11_22, in_data_to_next_pe_11_23, 
                        in_data_to_next_pe_11_24, in_data_to_next_pe_11_25, in_data_to_next_pe_11_26, in_data_to_next_pe_11_27, 
                        in_data_to_next_pe_11_28, in_data_to_next_pe_11_29, in_data_to_next_pe_11_30, in_data_to_next_pe_11_31, 
                        
                        
                        in_data_to_next_pe_12_0, in_data_to_next_pe_12_1, in_data_to_next_pe_12_2, in_data_to_next_pe_12_3,  
                        in_data_to_next_pe_12_4, in_data_to_next_pe_12_5, in_data_to_next_pe_12_6, in_data_to_next_pe_12_7,
                        in_data_to_next_pe_12_8, in_data_to_next_pe_12_9, in_data_to_next_pe_12_10, in_data_to_next_pe_12_11,
                        in_data_to_next_pe_12_12, in_data_to_next_pe_12_13, in_data_to_next_pe_12_14, in_data_to_next_pe_12_15,
                        in_data_to_next_pe_12_16, in_data_to_next_pe_12_17, in_data_to_next_pe_12_18, in_data_to_next_pe_12_19, 
                        in_data_to_next_pe_12_20, in_data_to_next_pe_12_21, in_data_to_next_pe_12_22, in_data_to_next_pe_12_23, 
                        in_data_to_next_pe_12_24, in_data_to_next_pe_12_25, in_data_to_next_pe_12_26, in_data_to_next_pe_12_27, 
                        in_data_to_next_pe_12_28, in_data_to_next_pe_12_29, in_data_to_next_pe_12_30, in_data_to_next_pe_12_31, 
                        
                        
                        in_data_to_next_pe_13_0, in_data_to_next_pe_13_1, in_data_to_next_pe_13_2, in_data_to_next_pe_13_3,  
                        in_data_to_next_pe_13_4, in_data_to_next_pe_13_5, in_data_to_next_pe_13_6, in_data_to_next_pe_13_7,
                        in_data_to_next_pe_13_8, in_data_to_next_pe_13_9, in_data_to_next_pe_13_10, in_data_to_next_pe_13_11,
                        in_data_to_next_pe_13_12, in_data_to_next_pe_13_13, in_data_to_next_pe_13_14, in_data_to_next_pe_13_15,
                        in_data_to_next_pe_13_16, in_data_to_next_pe_13_17, in_data_to_next_pe_13_18, in_data_to_next_pe_13_19, 
                        in_data_to_next_pe_13_20, in_data_to_next_pe_13_21, in_data_to_next_pe_13_22, in_data_to_next_pe_13_23, 
                        in_data_to_next_pe_13_24, in_data_to_next_pe_13_25, in_data_to_next_pe_13_26, in_data_to_next_pe_13_27, 
                        in_data_to_next_pe_13_28, in_data_to_next_pe_13_29, in_data_to_next_pe_13_30, in_data_to_next_pe_13_31, 
                        
                        
                        in_data_to_next_pe_14_0, in_data_to_next_pe_14_1, in_data_to_next_pe_14_2, in_data_to_next_pe_14_3,  
                        in_data_to_next_pe_14_4, in_data_to_next_pe_14_5, in_data_to_next_pe_14_6, in_data_to_next_pe_14_7,
                        in_data_to_next_pe_14_8, in_data_to_next_pe_14_9, in_data_to_next_pe_14_10, in_data_to_next_pe_14_11,
                        in_data_to_next_pe_14_12, in_data_to_next_pe_14_13, in_data_to_next_pe_14_14, in_data_to_next_pe_14_15,
                        in_data_to_next_pe_14_16, in_data_to_next_pe_14_17, in_data_to_next_pe_14_18, in_data_to_next_pe_14_19, 
                        in_data_to_next_pe_14_20, in_data_to_next_pe_14_21, in_data_to_next_pe_14_22, in_data_to_next_pe_14_23, 
                        in_data_to_next_pe_14_24, in_data_to_next_pe_14_25, in_data_to_next_pe_14_26, in_data_to_next_pe_14_27, 
                        in_data_to_next_pe_14_28, in_data_to_next_pe_14_29, in_data_to_next_pe_14_30, in_data_to_next_pe_14_31, 
                        
                        
                        in_data_to_next_pe_15_0, in_data_to_next_pe_15_1, in_data_to_next_pe_15_2, in_data_to_next_pe_15_3,  
                        in_data_to_next_pe_15_4, in_data_to_next_pe_15_5, in_data_to_next_pe_15_6, in_data_to_next_pe_15_7,
                        in_data_to_next_pe_15_8, in_data_to_next_pe_15_9, in_data_to_next_pe_15_10, in_data_to_next_pe_15_11,
                        in_data_to_next_pe_15_12, in_data_to_next_pe_15_13, in_data_to_next_pe_15_14, in_data_to_next_pe_15_15,
                        in_data_to_next_pe_15_16, in_data_to_next_pe_15_17, in_data_to_next_pe_15_18, in_data_to_next_pe_15_19, 
                        in_data_to_next_pe_15_20, in_data_to_next_pe_15_21, in_data_to_next_pe_15_22, in_data_to_next_pe_15_23, 
                        in_data_to_next_pe_15_24, in_data_to_next_pe_15_25, in_data_to_next_pe_15_26, in_data_to_next_pe_15_27, 
                        in_data_to_next_pe_15_28, in_data_to_next_pe_15_29, in_data_to_next_pe_15_30, in_data_to_next_pe_15_31, 
                        
                        
                        in_data_to_next_pe_16_0, in_data_to_next_pe_16_1, in_data_to_next_pe_16_2, in_data_to_next_pe_16_3,  
                        in_data_to_next_pe_16_4, in_data_to_next_pe_16_5, in_data_to_next_pe_16_6, in_data_to_next_pe_16_7,
                        in_data_to_next_pe_16_8, in_data_to_next_pe_16_9, in_data_to_next_pe_16_10, in_data_to_next_pe_16_11,
                        in_data_to_next_pe_16_12, in_data_to_next_pe_16_13, in_data_to_next_pe_16_14, in_data_to_next_pe_16_15,
                        in_data_to_next_pe_16_16, in_data_to_next_pe_16_17, in_data_to_next_pe_16_18, in_data_to_next_pe_16_19, 
                        in_data_to_next_pe_16_20, in_data_to_next_pe_16_21, in_data_to_next_pe_16_22, in_data_to_next_pe_16_23, 
                        in_data_to_next_pe_16_24, in_data_to_next_pe_16_25, in_data_to_next_pe_16_26, in_data_to_next_pe_16_27, 
                        in_data_to_next_pe_16_28, in_data_to_next_pe_16_29, in_data_to_next_pe_16_30, in_data_to_next_pe_16_31, 
                        
                        
                        in_data_to_next_pe_17_0, in_data_to_next_pe_17_1, in_data_to_next_pe_17_2, in_data_to_next_pe_17_3,  
                        in_data_to_next_pe_17_4, in_data_to_next_pe_17_5, in_data_to_next_pe_17_6, in_data_to_next_pe_17_7,
                        in_data_to_next_pe_17_8, in_data_to_next_pe_17_9, in_data_to_next_pe_17_10, in_data_to_next_pe_17_11,
                        in_data_to_next_pe_17_12, in_data_to_next_pe_17_13, in_data_to_next_pe_17_14, in_data_to_next_pe_17_15,
                        in_data_to_next_pe_17_16, in_data_to_next_pe_17_17, in_data_to_next_pe_17_18, in_data_to_next_pe_17_19, 
                        in_data_to_next_pe_17_20, in_data_to_next_pe_17_21, in_data_to_next_pe_17_22, in_data_to_next_pe_17_23, 
                        in_data_to_next_pe_17_24, in_data_to_next_pe_17_25, in_data_to_next_pe_17_26, in_data_to_next_pe_17_27, 
                        in_data_to_next_pe_17_28, in_data_to_next_pe_17_29, in_data_to_next_pe_17_30, in_data_to_next_pe_17_31, 
                        
                        
                        in_data_to_next_pe_18_0, in_data_to_next_pe_18_1, in_data_to_next_pe_18_2, in_data_to_next_pe_18_3,  
                        in_data_to_next_pe_18_4, in_data_to_next_pe_18_5, in_data_to_next_pe_18_6, in_data_to_next_pe_18_7,
                        in_data_to_next_pe_18_8, in_data_to_next_pe_18_9, in_data_to_next_pe_18_10, in_data_to_next_pe_18_11,
                        in_data_to_next_pe_18_12, in_data_to_next_pe_18_13, in_data_to_next_pe_18_14, in_data_to_next_pe_18_15,
                        in_data_to_next_pe_18_16, in_data_to_next_pe_18_17, in_data_to_next_pe_18_18, in_data_to_next_pe_18_19, 
                        in_data_to_next_pe_18_20, in_data_to_next_pe_18_21, in_data_to_next_pe_18_22, in_data_to_next_pe_18_23, 
                        in_data_to_next_pe_18_24, in_data_to_next_pe_18_25, in_data_to_next_pe_18_26, in_data_to_next_pe_18_27, 
                        in_data_to_next_pe_18_28, in_data_to_next_pe_18_29, in_data_to_next_pe_18_30, in_data_to_next_pe_18_31, 
                        
                        
                        in_data_to_next_pe_19_0, in_data_to_next_pe_19_1, in_data_to_next_pe_19_2, in_data_to_next_pe_19_3,  
                        in_data_to_next_pe_19_4, in_data_to_next_pe_19_5, in_data_to_next_pe_19_6, in_data_to_next_pe_19_7,
                        in_data_to_next_pe_19_8, in_data_to_next_pe_19_9, in_data_to_next_pe_19_10, in_data_to_next_pe_19_11,
                        in_data_to_next_pe_19_12, in_data_to_next_pe_19_13, in_data_to_next_pe_19_14, in_data_to_next_pe_19_15,
                        in_data_to_next_pe_19_16, in_data_to_next_pe_19_17, in_data_to_next_pe_19_18, in_data_to_next_pe_19_19, 
                        in_data_to_next_pe_19_20, in_data_to_next_pe_19_21, in_data_to_next_pe_19_22, in_data_to_next_pe_19_23, 
                        in_data_to_next_pe_19_24, in_data_to_next_pe_19_25, in_data_to_next_pe_19_26, in_data_to_next_pe_19_27, 
                        in_data_to_next_pe_19_28, in_data_to_next_pe_19_29, in_data_to_next_pe_19_30, in_data_to_next_pe_19_31, 
                        
                        
                        in_data_to_next_pe_20_0, in_data_to_next_pe_20_1, in_data_to_next_pe_20_2, in_data_to_next_pe_20_3,  
                        in_data_to_next_pe_20_4, in_data_to_next_pe_20_5, in_data_to_next_pe_20_6, in_data_to_next_pe_20_7,
                        in_data_to_next_pe_20_8, in_data_to_next_pe_20_9, in_data_to_next_pe_20_10, in_data_to_next_pe_20_11,
                        in_data_to_next_pe_20_12, in_data_to_next_pe_20_13, in_data_to_next_pe_20_14, in_data_to_next_pe_20_15,
                        in_data_to_next_pe_20_16, in_data_to_next_pe_20_17, in_data_to_next_pe_20_18, in_data_to_next_pe_20_19, 
                        in_data_to_next_pe_20_20, in_data_to_next_pe_20_21, in_data_to_next_pe_20_22, in_data_to_next_pe_20_23, 
                        in_data_to_next_pe_20_24, in_data_to_next_pe_20_25, in_data_to_next_pe_20_26, in_data_to_next_pe_20_27, 
                        in_data_to_next_pe_20_28, in_data_to_next_pe_20_29, in_data_to_next_pe_20_30, in_data_to_next_pe_20_31, 
                        
                        
                        in_data_to_next_pe_21_0, in_data_to_next_pe_21_1, in_data_to_next_pe_21_2, in_data_to_next_pe_21_3,  
                        in_data_to_next_pe_21_4, in_data_to_next_pe_21_5, in_data_to_next_pe_21_6, in_data_to_next_pe_21_7,
                        in_data_to_next_pe_21_8, in_data_to_next_pe_21_9, in_data_to_next_pe_21_10, in_data_to_next_pe_21_11,
                        in_data_to_next_pe_21_12, in_data_to_next_pe_21_13, in_data_to_next_pe_21_14, in_data_to_next_pe_21_15,
                        in_data_to_next_pe_21_16, in_data_to_next_pe_21_17, in_data_to_next_pe_21_18, in_data_to_next_pe_21_19, 
                        in_data_to_next_pe_21_20, in_data_to_next_pe_21_21, in_data_to_next_pe_21_22, in_data_to_next_pe_21_23, 
                        in_data_to_next_pe_21_24, in_data_to_next_pe_21_25, in_data_to_next_pe_21_26, in_data_to_next_pe_21_27, 
                        in_data_to_next_pe_21_28, in_data_to_next_pe_21_29, in_data_to_next_pe_21_30, in_data_to_next_pe_21_31, 
                        
                        
                        in_data_to_next_pe_22_0, in_data_to_next_pe_22_1, in_data_to_next_pe_22_2, in_data_to_next_pe_22_3,  
                        in_data_to_next_pe_22_4, in_data_to_next_pe_22_5, in_data_to_next_pe_22_6, in_data_to_next_pe_22_7,
                        in_data_to_next_pe_22_8, in_data_to_next_pe_22_9, in_data_to_next_pe_22_10, in_data_to_next_pe_22_11,
                        in_data_to_next_pe_22_12, in_data_to_next_pe_22_13, in_data_to_next_pe_22_14, in_data_to_next_pe_22_15,
                        in_data_to_next_pe_22_16, in_data_to_next_pe_22_17, in_data_to_next_pe_22_18, in_data_to_next_pe_22_19, 
                        in_data_to_next_pe_22_20, in_data_to_next_pe_22_21, in_data_to_next_pe_22_22, in_data_to_next_pe_22_23, 
                        in_data_to_next_pe_22_24, in_data_to_next_pe_22_25, in_data_to_next_pe_22_26, in_data_to_next_pe_22_27, 
                        in_data_to_next_pe_22_28, in_data_to_next_pe_22_29, in_data_to_next_pe_22_30, in_data_to_next_pe_22_31, 
                        
                        
                        in_data_to_next_pe_23_0, in_data_to_next_pe_23_1, in_data_to_next_pe_23_2, in_data_to_next_pe_23_3,  
                        in_data_to_next_pe_23_4, in_data_to_next_pe_23_5, in_data_to_next_pe_23_6, in_data_to_next_pe_23_7,
                        in_data_to_next_pe_23_8, in_data_to_next_pe_23_9, in_data_to_next_pe_23_10, in_data_to_next_pe_23_11,
                        in_data_to_next_pe_23_12, in_data_to_next_pe_23_13, in_data_to_next_pe_23_14, in_data_to_next_pe_23_15,
                        in_data_to_next_pe_23_16, in_data_to_next_pe_23_17, in_data_to_next_pe_23_18, in_data_to_next_pe_23_19, 
                        in_data_to_next_pe_23_20, in_data_to_next_pe_23_21, in_data_to_next_pe_23_22, in_data_to_next_pe_23_23, 
                        in_data_to_next_pe_23_24, in_data_to_next_pe_23_25, in_data_to_next_pe_23_26, in_data_to_next_pe_23_27, 
                        in_data_to_next_pe_23_28, in_data_to_next_pe_23_29, in_data_to_next_pe_23_30, in_data_to_next_pe_23_31, 
                        
                        
                        in_data_to_next_pe_24_0, in_data_to_next_pe_24_1, in_data_to_next_pe_24_2, in_data_to_next_pe_24_3,  
                        in_data_to_next_pe_24_4, in_data_to_next_pe_24_5, in_data_to_next_pe_24_6, in_data_to_next_pe_24_7,
                        in_data_to_next_pe_24_8, in_data_to_next_pe_24_9, in_data_to_next_pe_24_10, in_data_to_next_pe_24_11,
                        in_data_to_next_pe_24_12, in_data_to_next_pe_24_13, in_data_to_next_pe_24_14, in_data_to_next_pe_24_15,
                        in_data_to_next_pe_24_16, in_data_to_next_pe_24_17, in_data_to_next_pe_24_18, in_data_to_next_pe_24_19, 
                        in_data_to_next_pe_24_20, in_data_to_next_pe_24_21, in_data_to_next_pe_24_22, in_data_to_next_pe_24_23, 
                        in_data_to_next_pe_24_24, in_data_to_next_pe_24_25, in_data_to_next_pe_24_26, in_data_to_next_pe_24_27, 
                        in_data_to_next_pe_24_28, in_data_to_next_pe_24_29, in_data_to_next_pe_24_30, in_data_to_next_pe_24_31, 
                        
                        
                        in_data_to_next_pe_25_0, in_data_to_next_pe_25_1, in_data_to_next_pe_25_2, in_data_to_next_pe_25_3,  
                        in_data_to_next_pe_25_4, in_data_to_next_pe_25_5, in_data_to_next_pe_25_6, in_data_to_next_pe_25_7,
                        in_data_to_next_pe_25_8, in_data_to_next_pe_25_9, in_data_to_next_pe_25_10, in_data_to_next_pe_25_11,
                        in_data_to_next_pe_25_12, in_data_to_next_pe_25_13, in_data_to_next_pe_25_14, in_data_to_next_pe_25_15,
                        in_data_to_next_pe_25_16, in_data_to_next_pe_25_17, in_data_to_next_pe_25_18, in_data_to_next_pe_25_19, 
                        in_data_to_next_pe_25_20, in_data_to_next_pe_25_21, in_data_to_next_pe_25_22, in_data_to_next_pe_25_23, 
                        in_data_to_next_pe_25_24, in_data_to_next_pe_25_25, in_data_to_next_pe_25_26, in_data_to_next_pe_25_27, 
                        in_data_to_next_pe_25_28, in_data_to_next_pe_25_29, in_data_to_next_pe_25_30, in_data_to_next_pe_25_31, 
                        
                        
                        in_data_to_next_pe_26_0, in_data_to_next_pe_26_1, in_data_to_next_pe_26_2, in_data_to_next_pe_26_3,  
                        in_data_to_next_pe_26_4, in_data_to_next_pe_26_5, in_data_to_next_pe_26_6, in_data_to_next_pe_26_7,
                        in_data_to_next_pe_26_8, in_data_to_next_pe_26_9, in_data_to_next_pe_26_10, in_data_to_next_pe_26_11,
                        in_data_to_next_pe_26_12, in_data_to_next_pe_26_13, in_data_to_next_pe_26_14, in_data_to_next_pe_26_15,
                        in_data_to_next_pe_26_16, in_data_to_next_pe_26_17, in_data_to_next_pe_26_18, in_data_to_next_pe_26_19, 
                        in_data_to_next_pe_26_20, in_data_to_next_pe_26_21, in_data_to_next_pe_26_22, in_data_to_next_pe_26_23, 
                        in_data_to_next_pe_26_24, in_data_to_next_pe_26_25, in_data_to_next_pe_26_26, in_data_to_next_pe_26_27, 
                        in_data_to_next_pe_26_28, in_data_to_next_pe_26_29, in_data_to_next_pe_26_30, in_data_to_next_pe_26_31, 
                        
                        
                        in_data_to_next_pe_27_0, in_data_to_next_pe_27_1, in_data_to_next_pe_27_2, in_data_to_next_pe_27_3,  
                        in_data_to_next_pe_27_4, in_data_to_next_pe_27_5, in_data_to_next_pe_27_6, in_data_to_next_pe_27_7,
                        in_data_to_next_pe_27_8, in_data_to_next_pe_27_9, in_data_to_next_pe_27_10, in_data_to_next_pe_27_11,
                        in_data_to_next_pe_27_12, in_data_to_next_pe_27_13, in_data_to_next_pe_27_14, in_data_to_next_pe_27_15,
                        in_data_to_next_pe_27_16, in_data_to_next_pe_27_17, in_data_to_next_pe_27_18, in_data_to_next_pe_27_19, 
                        in_data_to_next_pe_27_20, in_data_to_next_pe_27_21, in_data_to_next_pe_27_22, in_data_to_next_pe_27_23, 
                        in_data_to_next_pe_27_24, in_data_to_next_pe_27_25, in_data_to_next_pe_27_26, in_data_to_next_pe_27_27, 
                        in_data_to_next_pe_27_28, in_data_to_next_pe_27_29, in_data_to_next_pe_27_30, in_data_to_next_pe_27_31, 
                        
                        
                        in_data_to_next_pe_28_0, in_data_to_next_pe_28_1, in_data_to_next_pe_28_2, in_data_to_next_pe_28_3,  
                        in_data_to_next_pe_28_4, in_data_to_next_pe_28_5, in_data_to_next_pe_28_6, in_data_to_next_pe_28_7,
                        in_data_to_next_pe_28_8, in_data_to_next_pe_28_9, in_data_to_next_pe_28_10, in_data_to_next_pe_28_11,
                        in_data_to_next_pe_28_12, in_data_to_next_pe_28_13, in_data_to_next_pe_28_14, in_data_to_next_pe_28_15,
                        in_data_to_next_pe_28_16, in_data_to_next_pe_28_17, in_data_to_next_pe_28_18, in_data_to_next_pe_28_19, 
                        in_data_to_next_pe_28_20, in_data_to_next_pe_28_21, in_data_to_next_pe_28_22, in_data_to_next_pe_28_23, 
                        in_data_to_next_pe_28_24, in_data_to_next_pe_28_25, in_data_to_next_pe_28_26, in_data_to_next_pe_28_27, 
                        in_data_to_next_pe_28_28, in_data_to_next_pe_28_29, in_data_to_next_pe_28_30, in_data_to_next_pe_28_31, 
                        
                        
                        in_data_to_next_pe_29_0, in_data_to_next_pe_29_1, in_data_to_next_pe_29_2, in_data_to_next_pe_29_3,  
                        in_data_to_next_pe_29_4, in_data_to_next_pe_29_5, in_data_to_next_pe_29_6, in_data_to_next_pe_29_7,
                        in_data_to_next_pe_29_8, in_data_to_next_pe_29_9, in_data_to_next_pe_29_10, in_data_to_next_pe_29_11,
                        in_data_to_next_pe_29_12, in_data_to_next_pe_29_13, in_data_to_next_pe_29_14, in_data_to_next_pe_29_15,
                        in_data_to_next_pe_29_16, in_data_to_next_pe_29_17, in_data_to_next_pe_29_18, in_data_to_next_pe_29_19, 
                        in_data_to_next_pe_29_20, in_data_to_next_pe_29_21, in_data_to_next_pe_29_22, in_data_to_next_pe_29_23, 
                        in_data_to_next_pe_29_24, in_data_to_next_pe_29_25, in_data_to_next_pe_29_26, in_data_to_next_pe_29_27, 
                        in_data_to_next_pe_29_28, in_data_to_next_pe_29_29, in_data_to_next_pe_29_30, in_data_to_next_pe_29_31, 
                        
                        
                        in_data_to_next_pe_30_0, in_data_to_next_pe_30_1, in_data_to_next_pe_30_2, in_data_to_next_pe_30_3,  
                        in_data_to_next_pe_30_4, in_data_to_next_pe_30_5, in_data_to_next_pe_30_6, in_data_to_next_pe_30_7,
                        in_data_to_next_pe_30_8, in_data_to_next_pe_30_9, in_data_to_next_pe_30_10, in_data_to_next_pe_30_11,
                        in_data_to_next_pe_30_12, in_data_to_next_pe_30_13, in_data_to_next_pe_30_14, in_data_to_next_pe_30_15,
                        in_data_to_next_pe_30_16, in_data_to_next_pe_30_17, in_data_to_next_pe_30_18, in_data_to_next_pe_30_19, 
                        in_data_to_next_pe_30_20, in_data_to_next_pe_30_21, in_data_to_next_pe_30_22, in_data_to_next_pe_30_23, 
                        in_data_to_next_pe_30_24, in_data_to_next_pe_30_25, in_data_to_next_pe_30_26, in_data_to_next_pe_30_27, 
                        in_data_to_next_pe_30_28, in_data_to_next_pe_30_29, in_data_to_next_pe_30_30, in_data_to_next_pe_30_31, 
                        
                        
                        in_data_to_next_pe_31_0, in_data_to_next_pe_31_1, in_data_to_next_pe_31_2, in_data_to_next_pe_31_3,  
                        in_data_to_next_pe_31_4, in_data_to_next_pe_31_5, in_data_to_next_pe_31_6, in_data_to_next_pe_31_7,
                        in_data_to_next_pe_31_8, in_data_to_next_pe_31_9, in_data_to_next_pe_31_10, in_data_to_next_pe_31_11,
                        in_data_to_next_pe_31_12, in_data_to_next_pe_31_13, in_data_to_next_pe_31_14, in_data_to_next_pe_31_15,
                        in_data_to_next_pe_31_16, in_data_to_next_pe_31_17, in_data_to_next_pe_31_18, in_data_to_next_pe_31_19, 
                        in_data_to_next_pe_31_20, in_data_to_next_pe_31_21, in_data_to_next_pe_31_22, in_data_to_next_pe_31_23, 
                        in_data_to_next_pe_31_24, in_data_to_next_pe_31_25, in_data_to_next_pe_31_26, in_data_to_next_pe_31_27, 
                        in_data_to_next_pe_31_28, in_data_to_next_pe_31_29, in_data_to_next_pe_31_30, in_data_to_next_pe_31_31,
                        
                        
        in_data_to_next_pe_32_0, in_data_to_next_pe_32_1, in_data_to_next_pe_32_2, in_data_to_next_pe_32_3,  
        in_data_to_next_pe_32_4, in_data_to_next_pe_32_5, in_data_to_next_pe_32_6, in_data_to_next_pe_32_7,
        in_data_to_next_pe_32_8, in_data_to_next_pe_32_9, in_data_to_next_pe_32_10, in_data_to_next_pe_32_11,
        in_data_to_next_pe_32_12, in_data_to_next_pe_32_13, in_data_to_next_pe_32_14, in_data_to_next_pe_32_15,
        in_data_to_next_pe_32_16, in_data_to_next_pe_32_17, in_data_to_next_pe_32_18, in_data_to_next_pe_32_19, 
        in_data_to_next_pe_32_20, in_data_to_next_pe_32_21, in_data_to_next_pe_32_22, in_data_to_next_pe_32_23, 
        in_data_to_next_pe_32_24, in_data_to_next_pe_32_25, in_data_to_next_pe_32_26, in_data_to_next_pe_32_27, 
        in_data_to_next_pe_32_28, in_data_to_next_pe_32_29, in_data_to_next_pe_32_30, in_data_to_next_pe_32_31,
        
        in_data_to_next_pe_33_0, in_data_to_next_pe_33_1, in_data_to_next_pe_33_2, in_data_to_next_pe_33_3,  
        in_data_to_next_pe_33_4, in_data_to_next_pe_33_5, in_data_to_next_pe_33_6, in_data_to_next_pe_33_7,
        in_data_to_next_pe_33_8, in_data_to_next_pe_33_9, in_data_to_next_pe_33_10, in_data_to_next_pe_33_11,
        in_data_to_next_pe_33_12, in_data_to_next_pe_33_13, in_data_to_next_pe_33_14, in_data_to_next_pe_33_15,
        in_data_to_next_pe_33_16, in_data_to_next_pe_33_17, in_data_to_next_pe_33_18, in_data_to_next_pe_33_19, 
        in_data_to_next_pe_33_20, in_data_to_next_pe_33_21, in_data_to_next_pe_33_22, in_data_to_next_pe_33_23, 
        in_data_to_next_pe_33_24, in_data_to_next_pe_33_25, in_data_to_next_pe_33_26, in_data_to_next_pe_33_27, 
        in_data_to_next_pe_33_28, in_data_to_next_pe_33_29, in_data_to_next_pe_33_30, in_data_to_next_pe_33_31,
        
        in_data_to_next_pe_34_0, in_data_to_next_pe_34_1, in_data_to_next_pe_34_2, in_data_to_next_pe_34_3,  
        in_data_to_next_pe_34_4, in_data_to_next_pe_34_5, in_data_to_next_pe_34_6, in_data_to_next_pe_34_7,
        in_data_to_next_pe_34_8, in_data_to_next_pe_34_9, in_data_to_next_pe_34_10, in_data_to_next_pe_34_11,
        in_data_to_next_pe_34_12, in_data_to_next_pe_34_13, in_data_to_next_pe_34_14, in_data_to_next_pe_34_15,
        in_data_to_next_pe_34_16, in_data_to_next_pe_34_17, in_data_to_next_pe_34_18, in_data_to_next_pe_34_19, 
        in_data_to_next_pe_34_20, in_data_to_next_pe_34_21, in_data_to_next_pe_34_22, in_data_to_next_pe_34_23, 
        in_data_to_next_pe_34_24, in_data_to_next_pe_34_25, in_data_to_next_pe_34_26, in_data_to_next_pe_34_27, 
        in_data_to_next_pe_34_28, in_data_to_next_pe_34_29, in_data_to_next_pe_34_30, in_data_to_next_pe_34_31,
        
        in_data_to_next_pe_35_0, in_data_to_next_pe_35_1, in_data_to_next_pe_35_2, in_data_to_next_pe_35_3,  
        in_data_to_next_pe_35_4, in_data_to_next_pe_35_5, in_data_to_next_pe_35_6, in_data_to_next_pe_35_7,
        in_data_to_next_pe_35_8, in_data_to_next_pe_35_9, in_data_to_next_pe_35_10, in_data_to_next_pe_35_11,
        in_data_to_next_pe_35_12, in_data_to_next_pe_35_13, in_data_to_next_pe_35_14, in_data_to_next_pe_35_15,
        in_data_to_next_pe_35_16, in_data_to_next_pe_35_17, in_data_to_next_pe_35_18, in_data_to_next_pe_35_19, 
        in_data_to_next_pe_35_20, in_data_to_next_pe_35_21, in_data_to_next_pe_35_22, in_data_to_next_pe_35_23, 
        in_data_to_next_pe_35_24, in_data_to_next_pe_35_25, in_data_to_next_pe_35_26, in_data_to_next_pe_35_27, 
        in_data_to_next_pe_35_28, in_data_to_next_pe_35_29, in_data_to_next_pe_35_30, in_data_to_next_pe_35_31,
        
        in_data_to_next_pe_36_0, in_data_to_next_pe_36_1, in_data_to_next_pe_36_2, in_data_to_next_pe_36_3,  
        in_data_to_next_pe_36_4, in_data_to_next_pe_36_5, in_data_to_next_pe_36_6, in_data_to_next_pe_36_7,
        in_data_to_next_pe_36_8, in_data_to_next_pe_36_9, in_data_to_next_pe_36_10, in_data_to_next_pe_36_11,
        in_data_to_next_pe_36_12, in_data_to_next_pe_36_13, in_data_to_next_pe_36_14, in_data_to_next_pe_36_15,
        in_data_to_next_pe_36_16, in_data_to_next_pe_36_17, in_data_to_next_pe_36_18, in_data_to_next_pe_36_19, 
        in_data_to_next_pe_36_20, in_data_to_next_pe_36_21, in_data_to_next_pe_36_22, in_data_to_next_pe_36_23, 
        in_data_to_next_pe_36_24, in_data_to_next_pe_36_25, in_data_to_next_pe_36_26, in_data_to_next_pe_36_27, 
        in_data_to_next_pe_36_28, in_data_to_next_pe_36_29, in_data_to_next_pe_36_30, in_data_to_next_pe_36_31,
        
        in_data_to_next_pe_37_0, in_data_to_next_pe_37_1, in_data_to_next_pe_37_2, in_data_to_next_pe_37_3,  
        in_data_to_next_pe_37_4, in_data_to_next_pe_37_5, in_data_to_next_pe_37_6, in_data_to_next_pe_37_7,
        in_data_to_next_pe_37_8, in_data_to_next_pe_37_9, in_data_to_next_pe_37_10, in_data_to_next_pe_37_11,
        in_data_to_next_pe_37_12, in_data_to_next_pe_37_13, in_data_to_next_pe_37_14, in_data_to_next_pe_37_15,
        in_data_to_next_pe_37_16, in_data_to_next_pe_37_17, in_data_to_next_pe_37_18, in_data_to_next_pe_37_19, 
        in_data_to_next_pe_37_20, in_data_to_next_pe_37_21, in_data_to_next_pe_37_22, in_data_to_next_pe_37_23, 
        in_data_to_next_pe_37_24, in_data_to_next_pe_37_25, in_data_to_next_pe_37_26, in_data_to_next_pe_37_27, 
        in_data_to_next_pe_37_28, in_data_to_next_pe_37_29, in_data_to_next_pe_37_30, in_data_to_next_pe_37_31,
        
        in_data_to_next_pe_38_0, in_data_to_next_pe_38_1, in_data_to_next_pe_38_2, in_data_to_next_pe_38_3,  
        in_data_to_next_pe_38_4, in_data_to_next_pe_38_5, in_data_to_next_pe_38_6, in_data_to_next_pe_38_7,
        in_data_to_next_pe_38_8, in_data_to_next_pe_38_9, in_data_to_next_pe_38_10, in_data_to_next_pe_38_11,
        in_data_to_next_pe_38_12, in_data_to_next_pe_38_13, in_data_to_next_pe_38_14, in_data_to_next_pe_38_15,
        in_data_to_next_pe_38_16, in_data_to_next_pe_38_17, in_data_to_next_pe_38_18, in_data_to_next_pe_38_19, 
        in_data_to_next_pe_38_20, in_data_to_next_pe_38_21, in_data_to_next_pe_38_22, in_data_to_next_pe_38_23, 
        in_data_to_next_pe_38_24, in_data_to_next_pe_38_25, in_data_to_next_pe_38_26, in_data_to_next_pe_38_27, 
        in_data_to_next_pe_38_28, in_data_to_next_pe_38_29, in_data_to_next_pe_38_30, in_data_to_next_pe_38_31,
        
        in_data_to_next_pe_39_0, in_data_to_next_pe_39_1, in_data_to_next_pe_39_2, in_data_to_next_pe_39_3,  
        in_data_to_next_pe_39_4, in_data_to_next_pe_39_5, in_data_to_next_pe_39_6, in_data_to_next_pe_39_7,
        in_data_to_next_pe_39_8, in_data_to_next_pe_39_9, in_data_to_next_pe_39_10, in_data_to_next_pe_39_11,
        in_data_to_next_pe_39_12, in_data_to_next_pe_39_13, in_data_to_next_pe_39_14, in_data_to_next_pe_39_15,
        in_data_to_next_pe_39_16, in_data_to_next_pe_39_17, in_data_to_next_pe_39_18, in_data_to_next_pe_39_19, 
        in_data_to_next_pe_39_20, in_data_to_next_pe_39_21, in_data_to_next_pe_39_22, in_data_to_next_pe_39_23, 
        in_data_to_next_pe_39_24, in_data_to_next_pe_39_25, in_data_to_next_pe_39_26, in_data_to_next_pe_39_27, 
        in_data_to_next_pe_39_28, in_data_to_next_pe_39_29, in_data_to_next_pe_39_30, in_data_to_next_pe_39_31,
        
        in_data_to_next_pe_40_0, in_data_to_next_pe_40_1, in_data_to_next_pe_40_2, in_data_to_next_pe_40_3,  
        in_data_to_next_pe_40_4, in_data_to_next_pe_40_5, in_data_to_next_pe_40_6, in_data_to_next_pe_40_7,
        in_data_to_next_pe_40_8, in_data_to_next_pe_40_9, in_data_to_next_pe_40_10, in_data_to_next_pe_40_11,
        in_data_to_next_pe_40_12, in_data_to_next_pe_40_13, in_data_to_next_pe_40_14, in_data_to_next_pe_40_15,
        in_data_to_next_pe_40_16, in_data_to_next_pe_40_17, in_data_to_next_pe_40_18, in_data_to_next_pe_40_19, 
        in_data_to_next_pe_40_20, in_data_to_next_pe_40_21, in_data_to_next_pe_40_22, in_data_to_next_pe_40_23, 
        in_data_to_next_pe_40_24, in_data_to_next_pe_40_25, in_data_to_next_pe_40_26, in_data_to_next_pe_40_27, 
        in_data_to_next_pe_40_28, in_data_to_next_pe_40_29, in_data_to_next_pe_40_30, in_data_to_next_pe_40_31,
        
        in_data_to_next_pe_41_0, in_data_to_next_pe_41_1, in_data_to_next_pe_41_2, in_data_to_next_pe_41_3,  
        in_data_to_next_pe_41_4, in_data_to_next_pe_41_5, in_data_to_next_pe_41_6, in_data_to_next_pe_41_7,
        in_data_to_next_pe_41_8, in_data_to_next_pe_41_9, in_data_to_next_pe_41_10, in_data_to_next_pe_41_11,
        in_data_to_next_pe_41_12, in_data_to_next_pe_41_13, in_data_to_next_pe_41_14, in_data_to_next_pe_41_15,
        in_data_to_next_pe_41_16, in_data_to_next_pe_41_17, in_data_to_next_pe_41_18, in_data_to_next_pe_41_19, 
        in_data_to_next_pe_41_20, in_data_to_next_pe_41_21, in_data_to_next_pe_41_22, in_data_to_next_pe_41_23, 
        in_data_to_next_pe_41_24, in_data_to_next_pe_41_25, in_data_to_next_pe_41_26, in_data_to_next_pe_41_27, 
        in_data_to_next_pe_41_28, in_data_to_next_pe_41_29, in_data_to_next_pe_41_30, in_data_to_next_pe_41_31,
        
        in_data_to_next_pe_42_0, in_data_to_next_pe_42_1, in_data_to_next_pe_42_2, in_data_to_next_pe_42_3,  
        in_data_to_next_pe_42_4, in_data_to_next_pe_42_5, in_data_to_next_pe_42_6, in_data_to_next_pe_42_7,
        in_data_to_next_pe_42_8, in_data_to_next_pe_42_9, in_data_to_next_pe_42_10, in_data_to_next_pe_42_11,
        in_data_to_next_pe_42_12, in_data_to_next_pe_42_13, in_data_to_next_pe_42_14, in_data_to_next_pe_42_15,
        in_data_to_next_pe_42_16, in_data_to_next_pe_42_17, in_data_to_next_pe_42_18, in_data_to_next_pe_42_19, 
        in_data_to_next_pe_42_20, in_data_to_next_pe_42_21, in_data_to_next_pe_42_22, in_data_to_next_pe_42_23, 
        in_data_to_next_pe_42_24, in_data_to_next_pe_42_25, in_data_to_next_pe_42_26, in_data_to_next_pe_42_27, 
        in_data_to_next_pe_42_28, in_data_to_next_pe_42_29, in_data_to_next_pe_42_30, in_data_to_next_pe_42_31,
        
        in_data_to_next_pe_43_0, in_data_to_next_pe_43_1, in_data_to_next_pe_43_2, in_data_to_next_pe_43_3,  
        in_data_to_next_pe_43_4, in_data_to_next_pe_43_5, in_data_to_next_pe_43_6, in_data_to_next_pe_43_7,
        in_data_to_next_pe_43_8, in_data_to_next_pe_43_9, in_data_to_next_pe_43_10, in_data_to_next_pe_43_11,
        in_data_to_next_pe_43_12, in_data_to_next_pe_43_13, in_data_to_next_pe_43_14, in_data_to_next_pe_43_15,
        in_data_to_next_pe_43_16, in_data_to_next_pe_43_17, in_data_to_next_pe_43_18, in_data_to_next_pe_43_19, 
        in_data_to_next_pe_43_20, in_data_to_next_pe_43_21, in_data_to_next_pe_43_22, in_data_to_next_pe_43_23, 
        in_data_to_next_pe_43_24, in_data_to_next_pe_43_25, in_data_to_next_pe_43_26, in_data_to_next_pe_43_27, 
        in_data_to_next_pe_43_28, in_data_to_next_pe_43_29, in_data_to_next_pe_43_30, in_data_to_next_pe_43_31,
        
        in_data_to_next_pe_44_0, in_data_to_next_pe_44_1, in_data_to_next_pe_44_2, in_data_to_next_pe_44_3,  
        in_data_to_next_pe_44_4, in_data_to_next_pe_44_5, in_data_to_next_pe_44_6, in_data_to_next_pe_44_7,
        in_data_to_next_pe_44_8, in_data_to_next_pe_44_9, in_data_to_next_pe_44_10, in_data_to_next_pe_44_11,
        in_data_to_next_pe_44_12, in_data_to_next_pe_44_13, in_data_to_next_pe_44_14, in_data_to_next_pe_44_15,
        in_data_to_next_pe_44_16, in_data_to_next_pe_44_17, in_data_to_next_pe_44_18, in_data_to_next_pe_44_19, 
        in_data_to_next_pe_44_20, in_data_to_next_pe_44_21, in_data_to_next_pe_44_22, in_data_to_next_pe_44_23, 
        in_data_to_next_pe_44_24, in_data_to_next_pe_44_25, in_data_to_next_pe_44_26, in_data_to_next_pe_44_27, 
        in_data_to_next_pe_44_28, in_data_to_next_pe_44_29, in_data_to_next_pe_44_30, in_data_to_next_pe_44_31,
        
        in_data_to_next_pe_45_0, in_data_to_next_pe_45_1, in_data_to_next_pe_45_2, in_data_to_next_pe_45_3,  
        in_data_to_next_pe_45_4, in_data_to_next_pe_45_5, in_data_to_next_pe_45_6, in_data_to_next_pe_45_7,
        in_data_to_next_pe_45_8, in_data_to_next_pe_45_9, in_data_to_next_pe_45_10, in_data_to_next_pe_45_11,
        in_data_to_next_pe_45_12, in_data_to_next_pe_45_13, in_data_to_next_pe_45_14, in_data_to_next_pe_45_15,
        in_data_to_next_pe_45_16, in_data_to_next_pe_45_17, in_data_to_next_pe_45_18, in_data_to_next_pe_45_19, 
        in_data_to_next_pe_45_20, in_data_to_next_pe_45_21, in_data_to_next_pe_45_22, in_data_to_next_pe_45_23, 
        in_data_to_next_pe_45_24, in_data_to_next_pe_45_25, in_data_to_next_pe_45_26, in_data_to_next_pe_45_27, 
        in_data_to_next_pe_45_28, in_data_to_next_pe_45_29, in_data_to_next_pe_45_30, in_data_to_next_pe_45_31,
        
        in_data_to_next_pe_46_0, in_data_to_next_pe_46_1, in_data_to_next_pe_46_2, in_data_to_next_pe_46_3,  
        in_data_to_next_pe_46_4, in_data_to_next_pe_46_5, in_data_to_next_pe_46_6, in_data_to_next_pe_46_7,
        in_data_to_next_pe_46_8, in_data_to_next_pe_46_9, in_data_to_next_pe_46_10, in_data_to_next_pe_46_11,
        in_data_to_next_pe_46_12, in_data_to_next_pe_46_13, in_data_to_next_pe_46_14, in_data_to_next_pe_46_15,
        in_data_to_next_pe_46_16, in_data_to_next_pe_46_17, in_data_to_next_pe_46_18, in_data_to_next_pe_46_19, 
        in_data_to_next_pe_46_20, in_data_to_next_pe_46_21, in_data_to_next_pe_46_22, in_data_to_next_pe_46_23, 
        in_data_to_next_pe_46_24, in_data_to_next_pe_46_25, in_data_to_next_pe_46_26, in_data_to_next_pe_46_27, 
        in_data_to_next_pe_46_28, in_data_to_next_pe_46_29, in_data_to_next_pe_46_30, in_data_to_next_pe_46_31,
        
        in_data_to_next_pe_47_0, in_data_to_next_pe_47_1, in_data_to_next_pe_47_2, in_data_to_next_pe_47_3,  
        in_data_to_next_pe_47_4, in_data_to_next_pe_47_5, in_data_to_next_pe_47_6, in_data_to_next_pe_47_7,
        in_data_to_next_pe_47_8, in_data_to_next_pe_47_9, in_data_to_next_pe_47_10, in_data_to_next_pe_47_11,
        in_data_to_next_pe_47_12, in_data_to_next_pe_47_13, in_data_to_next_pe_47_14, in_data_to_next_pe_47_15,
        in_data_to_next_pe_47_16, in_data_to_next_pe_47_17, in_data_to_next_pe_47_18, in_data_to_next_pe_47_19, 
        in_data_to_next_pe_47_20, in_data_to_next_pe_47_21, in_data_to_next_pe_47_22, in_data_to_next_pe_47_23, 
        in_data_to_next_pe_47_24, in_data_to_next_pe_47_25, in_data_to_next_pe_47_26, in_data_to_next_pe_47_27, 
        in_data_to_next_pe_47_28, in_data_to_next_pe_47_29, in_data_to_next_pe_47_30, in_data_to_next_pe_47_31,
        
        in_data_to_next_pe_48_0, in_data_to_next_pe_48_1, in_data_to_next_pe_48_2, in_data_to_next_pe_48_3,  
        in_data_to_next_pe_48_4, in_data_to_next_pe_48_5, in_data_to_next_pe_48_6, in_data_to_next_pe_48_7,
        in_data_to_next_pe_48_8, in_data_to_next_pe_48_9, in_data_to_next_pe_48_10, in_data_to_next_pe_48_11,
        in_data_to_next_pe_48_12, in_data_to_next_pe_48_13, in_data_to_next_pe_48_14, in_data_to_next_pe_48_15,
        in_data_to_next_pe_48_16, in_data_to_next_pe_48_17, in_data_to_next_pe_48_18, in_data_to_next_pe_48_19, 
        in_data_to_next_pe_48_20, in_data_to_next_pe_48_21, in_data_to_next_pe_48_22, in_data_to_next_pe_48_23, 
        in_data_to_next_pe_48_24, in_data_to_next_pe_48_25, in_data_to_next_pe_48_26, in_data_to_next_pe_48_27, 
        in_data_to_next_pe_48_28, in_data_to_next_pe_48_29, in_data_to_next_pe_48_30, in_data_to_next_pe_48_31,
        
        in_data_to_next_pe_49_0, in_data_to_next_pe_49_1, in_data_to_next_pe_49_2, in_data_to_next_pe_49_3,  
        in_data_to_next_pe_49_4, in_data_to_next_pe_49_5, in_data_to_next_pe_49_6, in_data_to_next_pe_49_7,
        in_data_to_next_pe_49_8, in_data_to_next_pe_49_9, in_data_to_next_pe_49_10, in_data_to_next_pe_49_11,
        in_data_to_next_pe_49_12, in_data_to_next_pe_49_13, in_data_to_next_pe_49_14, in_data_to_next_pe_49_15,
        in_data_to_next_pe_49_16, in_data_to_next_pe_49_17, in_data_to_next_pe_49_18, in_data_to_next_pe_49_19, 
        in_data_to_next_pe_49_20, in_data_to_next_pe_49_21, in_data_to_next_pe_49_22, in_data_to_next_pe_49_23, 
        in_data_to_next_pe_49_24, in_data_to_next_pe_49_25, in_data_to_next_pe_49_26, in_data_to_next_pe_49_27, 
        in_data_to_next_pe_49_28, in_data_to_next_pe_49_29, in_data_to_next_pe_49_30, in_data_to_next_pe_49_31,
        
        in_data_to_next_pe_50_0, in_data_to_next_pe_50_1, in_data_to_next_pe_50_2, in_data_to_next_pe_50_3,  
        in_data_to_next_pe_50_4, in_data_to_next_pe_50_5, in_data_to_next_pe_50_6, in_data_to_next_pe_50_7,
        in_data_to_next_pe_50_8, in_data_to_next_pe_50_9, in_data_to_next_pe_50_10, in_data_to_next_pe_50_11,
        in_data_to_next_pe_50_12, in_data_to_next_pe_50_13, in_data_to_next_pe_50_14, in_data_to_next_pe_50_15,
        in_data_to_next_pe_50_16, in_data_to_next_pe_50_17, in_data_to_next_pe_50_18, in_data_to_next_pe_50_19, 
        in_data_to_next_pe_50_20, in_data_to_next_pe_50_21, in_data_to_next_pe_50_22, in_data_to_next_pe_50_23, 
        in_data_to_next_pe_50_24, in_data_to_next_pe_50_25, in_data_to_next_pe_50_26, in_data_to_next_pe_50_27, 
        in_data_to_next_pe_50_28, in_data_to_next_pe_50_29, in_data_to_next_pe_50_30, in_data_to_next_pe_50_31,
        
        in_data_to_next_pe_51_0, in_data_to_next_pe_51_1, in_data_to_next_pe_51_2, in_data_to_next_pe_51_3,  
        in_data_to_next_pe_51_4, in_data_to_next_pe_51_5, in_data_to_next_pe_51_6, in_data_to_next_pe_51_7,
        in_data_to_next_pe_51_8, in_data_to_next_pe_51_9, in_data_to_next_pe_51_10, in_data_to_next_pe_51_11,
        in_data_to_next_pe_51_12, in_data_to_next_pe_51_13, in_data_to_next_pe_51_14, in_data_to_next_pe_51_15,
        in_data_to_next_pe_51_16, in_data_to_next_pe_51_17, in_data_to_next_pe_51_18, in_data_to_next_pe_51_19, 
        in_data_to_next_pe_51_20, in_data_to_next_pe_51_21, in_data_to_next_pe_51_22, in_data_to_next_pe_51_23, 
        in_data_to_next_pe_51_24, in_data_to_next_pe_51_25, in_data_to_next_pe_51_26, in_data_to_next_pe_51_27, 
        in_data_to_next_pe_51_28, in_data_to_next_pe_51_29, in_data_to_next_pe_51_30, in_data_to_next_pe_51_31,
        
        in_data_to_next_pe_52_0, in_data_to_next_pe_52_1, in_data_to_next_pe_52_2, in_data_to_next_pe_52_3,  
        in_data_to_next_pe_52_4, in_data_to_next_pe_52_5, in_data_to_next_pe_52_6, in_data_to_next_pe_52_7,
        in_data_to_next_pe_52_8, in_data_to_next_pe_52_9, in_data_to_next_pe_52_10, in_data_to_next_pe_52_11,
        in_data_to_next_pe_52_12, in_data_to_next_pe_52_13, in_data_to_next_pe_52_14, in_data_to_next_pe_52_15,
        in_data_to_next_pe_52_16, in_data_to_next_pe_52_17, in_data_to_next_pe_52_18, in_data_to_next_pe_52_19, 
        in_data_to_next_pe_52_20, in_data_to_next_pe_52_21, in_data_to_next_pe_52_22, in_data_to_next_pe_52_23, 
        in_data_to_next_pe_52_24, in_data_to_next_pe_52_25, in_data_to_next_pe_52_26, in_data_to_next_pe_52_27, 
        in_data_to_next_pe_52_28, in_data_to_next_pe_52_29, in_data_to_next_pe_52_30, in_data_to_next_pe_52_31,
        
        in_data_to_next_pe_53_0, in_data_to_next_pe_53_1, in_data_to_next_pe_53_2, in_data_to_next_pe_53_3,  
        in_data_to_next_pe_53_4, in_data_to_next_pe_53_5, in_data_to_next_pe_53_6, in_data_to_next_pe_53_7,
        in_data_to_next_pe_53_8, in_data_to_next_pe_53_9, in_data_to_next_pe_53_10, in_data_to_next_pe_53_11,
        in_data_to_next_pe_53_12, in_data_to_next_pe_53_13, in_data_to_next_pe_53_14, in_data_to_next_pe_53_15,
        in_data_to_next_pe_53_16, in_data_to_next_pe_53_17, in_data_to_next_pe_53_18, in_data_to_next_pe_53_19, 
        in_data_to_next_pe_53_20, in_data_to_next_pe_53_21, in_data_to_next_pe_53_22, in_data_to_next_pe_53_23, 
        in_data_to_next_pe_53_24, in_data_to_next_pe_53_25, in_data_to_next_pe_53_26, in_data_to_next_pe_53_27, 
        in_data_to_next_pe_53_28, in_data_to_next_pe_53_29, in_data_to_next_pe_53_30, in_data_to_next_pe_53_31,
        
        in_data_to_next_pe_54_0, in_data_to_next_pe_54_1, in_data_to_next_pe_54_2, in_data_to_next_pe_54_3,  
        in_data_to_next_pe_54_4, in_data_to_next_pe_54_5, in_data_to_next_pe_54_6, in_data_to_next_pe_54_7,
        in_data_to_next_pe_54_8, in_data_to_next_pe_54_9, in_data_to_next_pe_54_10, in_data_to_next_pe_54_11,
        in_data_to_next_pe_54_12, in_data_to_next_pe_54_13, in_data_to_next_pe_54_14, in_data_to_next_pe_54_15,
        in_data_to_next_pe_54_16, in_data_to_next_pe_54_17, in_data_to_next_pe_54_18, in_data_to_next_pe_54_19, 
        in_data_to_next_pe_54_20, in_data_to_next_pe_54_21, in_data_to_next_pe_54_22, in_data_to_next_pe_54_23, 
        in_data_to_next_pe_54_24, in_data_to_next_pe_54_25, in_data_to_next_pe_54_26, in_data_to_next_pe_54_27, 
        in_data_to_next_pe_54_28, in_data_to_next_pe_54_29, in_data_to_next_pe_54_30, in_data_to_next_pe_54_31,
        
        in_data_to_next_pe_55_0, in_data_to_next_pe_55_1, in_data_to_next_pe_55_2, in_data_to_next_pe_55_3,  
        in_data_to_next_pe_55_4, in_data_to_next_pe_55_5, in_data_to_next_pe_55_6, in_data_to_next_pe_55_7,
        in_data_to_next_pe_55_8, in_data_to_next_pe_55_9, in_data_to_next_pe_55_10, in_data_to_next_pe_55_11,
        in_data_to_next_pe_55_12, in_data_to_next_pe_55_13, in_data_to_next_pe_55_14, in_data_to_next_pe_55_15,
        in_data_to_next_pe_55_16, in_data_to_next_pe_55_17, in_data_to_next_pe_55_18, in_data_to_next_pe_55_19, 
        in_data_to_next_pe_55_20, in_data_to_next_pe_55_21, in_data_to_next_pe_55_22, in_data_to_next_pe_55_23, 
        in_data_to_next_pe_55_24, in_data_to_next_pe_55_25, in_data_to_next_pe_55_26, in_data_to_next_pe_55_27, 
        in_data_to_next_pe_55_28, in_data_to_next_pe_55_29, in_data_to_next_pe_55_30, in_data_to_next_pe_55_31,
        
        in_data_to_next_pe_56_0, in_data_to_next_pe_56_1, in_data_to_next_pe_56_2, in_data_to_next_pe_56_3,  
        in_data_to_next_pe_56_4, in_data_to_next_pe_56_5, in_data_to_next_pe_56_6, in_data_to_next_pe_56_7,
        in_data_to_next_pe_56_8, in_data_to_next_pe_56_9, in_data_to_next_pe_56_10, in_data_to_next_pe_56_11,
        in_data_to_next_pe_56_12, in_data_to_next_pe_56_13, in_data_to_next_pe_56_14, in_data_to_next_pe_56_15,
        in_data_to_next_pe_56_16, in_data_to_next_pe_56_17, in_data_to_next_pe_56_18, in_data_to_next_pe_56_19, 
        in_data_to_next_pe_56_20, in_data_to_next_pe_56_21, in_data_to_next_pe_56_22, in_data_to_next_pe_56_23, 
        in_data_to_next_pe_56_24, in_data_to_next_pe_56_25, in_data_to_next_pe_56_26, in_data_to_next_pe_56_27, 
        in_data_to_next_pe_56_28, in_data_to_next_pe_56_29, in_data_to_next_pe_56_30, in_data_to_next_pe_56_31,
        
        in_data_to_next_pe_57_0, in_data_to_next_pe_57_1, in_data_to_next_pe_57_2, in_data_to_next_pe_57_3,  
        in_data_to_next_pe_57_4, in_data_to_next_pe_57_5, in_data_to_next_pe_57_6, in_data_to_next_pe_57_7,
        in_data_to_next_pe_57_8, in_data_to_next_pe_57_9, in_data_to_next_pe_57_10, in_data_to_next_pe_57_11,
        in_data_to_next_pe_57_12, in_data_to_next_pe_57_13, in_data_to_next_pe_57_14, in_data_to_next_pe_57_15,
        in_data_to_next_pe_57_16, in_data_to_next_pe_57_17, in_data_to_next_pe_57_18, in_data_to_next_pe_57_19, 
        in_data_to_next_pe_57_20, in_data_to_next_pe_57_21, in_data_to_next_pe_57_22, in_data_to_next_pe_57_23, 
        in_data_to_next_pe_57_24, in_data_to_next_pe_57_25, in_data_to_next_pe_57_26, in_data_to_next_pe_57_27, 
        in_data_to_next_pe_57_28, in_data_to_next_pe_57_29, in_data_to_next_pe_57_30, in_data_to_next_pe_57_31,
        
        in_data_to_next_pe_58_0, in_data_to_next_pe_58_1, in_data_to_next_pe_58_2, in_data_to_next_pe_58_3,  
        in_data_to_next_pe_58_4, in_data_to_next_pe_58_5, in_data_to_next_pe_58_6, in_data_to_next_pe_58_7,
        in_data_to_next_pe_58_8, in_data_to_next_pe_58_9, in_data_to_next_pe_58_10, in_data_to_next_pe_58_11,
        in_data_to_next_pe_58_12, in_data_to_next_pe_58_13, in_data_to_next_pe_58_14, in_data_to_next_pe_58_15,
        in_data_to_next_pe_58_16, in_data_to_next_pe_58_17, in_data_to_next_pe_58_18, in_data_to_next_pe_58_19, 
        in_data_to_next_pe_58_20, in_data_to_next_pe_58_21, in_data_to_next_pe_58_22, in_data_to_next_pe_58_23, 
        in_data_to_next_pe_58_24, in_data_to_next_pe_58_25, in_data_to_next_pe_58_26, in_data_to_next_pe_58_27, 
        in_data_to_next_pe_58_28, in_data_to_next_pe_58_29, in_data_to_next_pe_58_30, in_data_to_next_pe_58_31,
        
        in_data_to_next_pe_59_0, in_data_to_next_pe_59_1, in_data_to_next_pe_59_2, in_data_to_next_pe_59_3,  
        in_data_to_next_pe_59_4, in_data_to_next_pe_59_5, in_data_to_next_pe_59_6, in_data_to_next_pe_59_7,
        in_data_to_next_pe_59_8, in_data_to_next_pe_59_9, in_data_to_next_pe_59_10, in_data_to_next_pe_59_11,
        in_data_to_next_pe_59_12, in_data_to_next_pe_59_13, in_data_to_next_pe_59_14, in_data_to_next_pe_59_15,
        in_data_to_next_pe_59_16, in_data_to_next_pe_59_17, in_data_to_next_pe_59_18, in_data_to_next_pe_59_19, 
        in_data_to_next_pe_59_20, in_data_to_next_pe_59_21, in_data_to_next_pe_59_22, in_data_to_next_pe_59_23, 
        in_data_to_next_pe_59_24, in_data_to_next_pe_59_25, in_data_to_next_pe_59_26, in_data_to_next_pe_59_27, 
        in_data_to_next_pe_59_28, in_data_to_next_pe_59_29, in_data_to_next_pe_59_30, in_data_to_next_pe_59_31,
        
        in_data_to_next_pe_60_0, in_data_to_next_pe_60_1, in_data_to_next_pe_60_2, in_data_to_next_pe_60_3,  
        in_data_to_next_pe_60_4, in_data_to_next_pe_60_5, in_data_to_next_pe_60_6, in_data_to_next_pe_60_7,
        in_data_to_next_pe_60_8, in_data_to_next_pe_60_9, in_data_to_next_pe_60_10, in_data_to_next_pe_60_11,
        in_data_to_next_pe_60_12, in_data_to_next_pe_60_13, in_data_to_next_pe_60_14, in_data_to_next_pe_60_15,
        in_data_to_next_pe_60_16, in_data_to_next_pe_60_17, in_data_to_next_pe_60_18, in_data_to_next_pe_60_19, 
        in_data_to_next_pe_60_20, in_data_to_next_pe_60_21, in_data_to_next_pe_60_22, in_data_to_next_pe_60_23, 
        in_data_to_next_pe_60_24, in_data_to_next_pe_60_25, in_data_to_next_pe_60_26, in_data_to_next_pe_60_27, 
        in_data_to_next_pe_60_28, in_data_to_next_pe_60_29, in_data_to_next_pe_60_30, in_data_to_next_pe_60_31,
        
        in_data_to_next_pe_61_0, in_data_to_next_pe_61_1, in_data_to_next_pe_61_2, in_data_to_next_pe_61_3,  
        in_data_to_next_pe_61_4, in_data_to_next_pe_61_5, in_data_to_next_pe_61_6, in_data_to_next_pe_61_7,
        in_data_to_next_pe_61_8, in_data_to_next_pe_61_9, in_data_to_next_pe_61_10, in_data_to_next_pe_61_11,
        in_data_to_next_pe_61_12, in_data_to_next_pe_61_13, in_data_to_next_pe_61_14, in_data_to_next_pe_61_15,
        in_data_to_next_pe_61_16, in_data_to_next_pe_61_17, in_data_to_next_pe_61_18, in_data_to_next_pe_61_19, 
        in_data_to_next_pe_61_20, in_data_to_next_pe_61_21, in_data_to_next_pe_61_22, in_data_to_next_pe_61_23, 
        in_data_to_next_pe_61_24, in_data_to_next_pe_61_25, in_data_to_next_pe_61_26, in_data_to_next_pe_61_27, 
        in_data_to_next_pe_61_28, in_data_to_next_pe_61_29, in_data_to_next_pe_61_30, in_data_to_next_pe_61_31,
        
        in_data_to_next_pe_62_0, in_data_to_next_pe_62_1, in_data_to_next_pe_62_2, in_data_to_next_pe_62_3,  
        in_data_to_next_pe_62_4, in_data_to_next_pe_62_5, in_data_to_next_pe_62_6, in_data_to_next_pe_62_7,
        in_data_to_next_pe_62_8, in_data_to_next_pe_62_9, in_data_to_next_pe_62_10, in_data_to_next_pe_62_11,
        in_data_to_next_pe_62_12, in_data_to_next_pe_62_13, in_data_to_next_pe_62_14, in_data_to_next_pe_62_15,
        in_data_to_next_pe_62_16, in_data_to_next_pe_62_17, in_data_to_next_pe_62_18, in_data_to_next_pe_62_19, 
        in_data_to_next_pe_62_20, in_data_to_next_pe_62_21, in_data_to_next_pe_62_22, in_data_to_next_pe_62_23, 
        in_data_to_next_pe_62_24, in_data_to_next_pe_62_25, in_data_to_next_pe_62_26, in_data_to_next_pe_62_27, 
        in_data_to_next_pe_62_28, in_data_to_next_pe_62_29, in_data_to_next_pe_62_30, in_data_to_next_pe_62_31,
        
        in_data_to_next_pe_63_0, in_data_to_next_pe_63_1, in_data_to_next_pe_63_2, in_data_to_next_pe_63_3,  
        in_data_to_next_pe_63_4, in_data_to_next_pe_63_5, in_data_to_next_pe_63_6, in_data_to_next_pe_63_7,
        in_data_to_next_pe_63_8, in_data_to_next_pe_63_9, in_data_to_next_pe_63_10, in_data_to_next_pe_63_11,
        in_data_to_next_pe_63_12, in_data_to_next_pe_63_13, in_data_to_next_pe_63_14, in_data_to_next_pe_63_15,
        in_data_to_next_pe_63_16, in_data_to_next_pe_63_17, in_data_to_next_pe_63_18, in_data_to_next_pe_63_19, 
        in_data_to_next_pe_63_20, in_data_to_next_pe_63_21, in_data_to_next_pe_63_22, in_data_to_next_pe_63_23, 
        in_data_to_next_pe_63_24, in_data_to_next_pe_63_25, in_data_to_next_pe_63_26, in_data_to_next_pe_63_27, 
        in_data_to_next_pe_63_28, in_data_to_next_pe_63_29, in_data_to_next_pe_63_30, in_data_to_next_pe_63_31;
        
        
        

wire                    row_1_en, row_2_en,  row_3_en,  row_4_en,  row_5_en,  row_6_en,  row_7_en, 
                        row_8_en, row_9_en, row_10_en, row_11_en, row_12_en, row_13_en, row_14_en, row_15_en,
                        row_16_en, row_17_en, row_18_en, row_19_en, row_20_en, row_21_en, row_22_en, row_23_en,
                        row_24_en, row_25_en, row_26_en, row_27_en, row_28_en, row_29_en, row_30_en, row_31_en,
                        row_32_en, row_33_en, row_34_en, row_35_en, row_36_en, row_37_en, row_38_en, row_39_en, 
                        row_40_en, row_41_en, row_42_en, row_43_en, row_44_en, row_45_en, row_46_en, row_47_en, 
                        row_48_en, row_49_en, row_50_en, row_51_en, row_52_en, row_53_en, row_54_en, row_55_en, 
                        row_56_en, row_57_en, row_58_en, row_59_en, row_60_en, row_61_en, row_62_en, row_63_en;
                        
PE_Row_B5   PE_R0_B5(   .clk(clk), .rst_n(rst_n), .new_weight_val(new_weight_val[0]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3), 
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11), 
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19), 
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23), 
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27), 
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31), 
                        .Slide_data_0(Slide_data_0), .Slide_data_1(Slide_data_1),
                        .Slide_data_2(Slide_data_2), .Slide_data_3(Slide_data_3), 
                        .Slide_data_4(Slide_data_4), .Slide_data_5(Slide_data_5),
                        .Slide_data_6(Slide_data_6), .Slide_data_7(Slide_data_7),
                        .Slide_data_8(Slide_data_8), .Slide_data_9(Slide_data_9),
                        .Slide_data_10(Slide_data_10), .Slide_data_11(Slide_data_11), 
                        .Slide_data_12(Slide_data_12), .Slide_data_13(Slide_data_13),
                        .Slide_data_14(Slide_data_14), .Slide_data_15(Slide_data_15),
                        .Slide_data_16(Slide_data_16), .Slide_data_17(Slide_data_17), 
                        .Slide_data_18(Slide_data_18), .Slide_data_19(Slide_data_19), 
                        .Slide_data_20(Slide_data_20), .Slide_data_21(Slide_data_21), 
                        .Slide_data_22(Slide_data_22), .Slide_data_23(Slide_data_23), 
                        .Slide_data_24(Slide_data_24), .Slide_data_25(Slide_data_25), 
                        .Slide_data_26(Slide_data_26), .Slide_data_27(Slide_data_27), 
                        .Slide_data_28(Slide_data_28), .Slide_data_29(Slide_data_29), 
                        .Slide_data_30(Slide_data_30), .Slide_data_31(Slide_data_31), 
                        .result(o_0),
                        .in_data_to_next_pe_0(in_data_to_next_pe_1_0), .in_data_to_next_pe_1(in_data_to_next_pe_1_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_1_2), .in_data_to_next_pe_3(in_data_to_next_pe_1_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_1_4), .in_data_to_next_pe_5(in_data_to_next_pe_1_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_1_6), .in_data_to_next_pe_7(in_data_to_next_pe_1_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_1_8), .in_data_to_next_pe_9(in_data_to_next_pe_1_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_1_10), .in_data_to_next_pe_11(in_data_to_next_pe_1_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_1_12), .in_data_to_next_pe_13(in_data_to_next_pe_1_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_1_14), .in_data_to_next_pe_15(in_data_to_next_pe_1_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_1_16), .in_data_to_next_pe_17(in_data_to_next_pe_1_17), 
                        .in_data_to_next_pe_18(in_data_to_next_pe_1_18), .in_data_to_next_pe_19(in_data_to_next_pe_1_19), 
                        .in_data_to_next_pe_20(in_data_to_next_pe_1_20), .in_data_to_next_pe_21(in_data_to_next_pe_1_21), 
                        .in_data_to_next_pe_22(in_data_to_next_pe_1_22), .in_data_to_next_pe_23(in_data_to_next_pe_1_23), 
                        .in_data_to_next_pe_24(in_data_to_next_pe_1_24), .in_data_to_next_pe_25(in_data_to_next_pe_1_25), 
                        .in_data_to_next_pe_26(in_data_to_next_pe_1_26), .in_data_to_next_pe_27(in_data_to_next_pe_1_27), 
                        .in_data_to_next_pe_28(in_data_to_next_pe_1_28), .in_data_to_next_pe_29(in_data_to_next_pe_1_29), 
                        .in_data_to_next_pe_30(in_data_to_next_pe_1_30), .in_data_to_next_pe_31(in_data_to_next_pe_1_31),
                        .next_row_en(row_1_en),  
                        .out_val(o_0_val)
);      

PE_Row_B5   PE_R1_B5(   .clk(clk), .rst_n(row_1_en), .new_weight_val(new_weight_val[1]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3), 
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11), 
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19), 
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23), 
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27), 
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31), 
                        .Slide_data_0(in_data_to_next_pe_1_0), .Slide_data_1(in_data_to_next_pe_1_1),
                        .Slide_data_2(in_data_to_next_pe_1_2), .Slide_data_3(in_data_to_next_pe_1_3), 
                        .Slide_data_4(in_data_to_next_pe_1_4), .Slide_data_5(in_data_to_next_pe_1_5),
                        .Slide_data_6(in_data_to_next_pe_1_6), .Slide_data_7(in_data_to_next_pe_1_7),
                        .Slide_data_8(in_data_to_next_pe_1_8), .Slide_data_9(in_data_to_next_pe_1_9),
                        .Slide_data_10(in_data_to_next_pe_1_10), .Slide_data_11(in_data_to_next_pe_1_11), 
                        .Slide_data_12(in_data_to_next_pe_1_12), .Slide_data_13(in_data_to_next_pe_1_13),
                        .Slide_data_14(in_data_to_next_pe_1_14), .Slide_data_15(in_data_to_next_pe_1_15),
                        .Slide_data_16(in_data_to_next_pe_1_16), .Slide_data_17(in_data_to_next_pe_1_17), 
                        .Slide_data_18(in_data_to_next_pe_1_18), .Slide_data_19(in_data_to_next_pe_1_19), 
                        .Slide_data_20(in_data_to_next_pe_1_20), .Slide_data_21(in_data_to_next_pe_1_21), 
                        .Slide_data_22(in_data_to_next_pe_1_22), .Slide_data_23(in_data_to_next_pe_1_23), 
                        .Slide_data_24(in_data_to_next_pe_1_24), .Slide_data_25(in_data_to_next_pe_1_25), 
                        .Slide_data_26(in_data_to_next_pe_1_26), .Slide_data_27(in_data_to_next_pe_1_27), 
                        .Slide_data_28(in_data_to_next_pe_1_28), .Slide_data_29(in_data_to_next_pe_1_29), 
                        .Slide_data_30(in_data_to_next_pe_1_30), .Slide_data_31(in_data_to_next_pe_1_31),
                        .result(o_1),
                        .in_data_to_next_pe_0(in_data_to_next_pe_2_0), .in_data_to_next_pe_1(in_data_to_next_pe_2_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_2_2), .in_data_to_next_pe_3(in_data_to_next_pe_2_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_2_4), .in_data_to_next_pe_5(in_data_to_next_pe_2_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_2_6), .in_data_to_next_pe_7(in_data_to_next_pe_2_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_2_8), .in_data_to_next_pe_9(in_data_to_next_pe_2_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_2_10), .in_data_to_next_pe_11(in_data_to_next_pe_2_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_2_12), .in_data_to_next_pe_13(in_data_to_next_pe_2_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_2_14), .in_data_to_next_pe_15(in_data_to_next_pe_2_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_2_16), .in_data_to_next_pe_17(in_data_to_next_pe_2_17), 
                        .in_data_to_next_pe_18(in_data_to_next_pe_2_18), .in_data_to_next_pe_19(in_data_to_next_pe_2_19), 
                        .in_data_to_next_pe_20(in_data_to_next_pe_2_20), .in_data_to_next_pe_21(in_data_to_next_pe_2_21), 
                        .in_data_to_next_pe_22(in_data_to_next_pe_2_22), .in_data_to_next_pe_23(in_data_to_next_pe_2_23), 
                        .in_data_to_next_pe_24(in_data_to_next_pe_2_24), .in_data_to_next_pe_25(in_data_to_next_pe_2_25), 
                        .in_data_to_next_pe_26(in_data_to_next_pe_2_26), .in_data_to_next_pe_27(in_data_to_next_pe_2_27), 
                        .in_data_to_next_pe_28(in_data_to_next_pe_2_28), .in_data_to_next_pe_29(in_data_to_next_pe_2_29), 
                        .in_data_to_next_pe_30(in_data_to_next_pe_2_30), .in_data_to_next_pe_31(in_data_to_next_pe_2_31), 
                        .next_row_en(row_2_en)
);

      
        PE_Row_B5   PE_R2_B5(   .clk(clk), .rst_n(row_2_en), .new_weight_val(new_weight_val[2]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_2_0), .Slide_data_1(in_data_to_next_pe_2_1),
                        .Slide_data_2(in_data_to_next_pe_2_2), .Slide_data_3(in_data_to_next_pe_2_3),
                        .Slide_data_4(in_data_to_next_pe_2_4), .Slide_data_5(in_data_to_next_pe_2_5),
                        .Slide_data_6(in_data_to_next_pe_2_6), .Slide_data_7(in_data_to_next_pe_2_7),
                        .Slide_data_8(in_data_to_next_pe_2_8), .Slide_data_9(in_data_to_next_pe_2_9),
                        .Slide_data_10(in_data_to_next_pe_2_10), .Slide_data_11(in_data_to_next_pe_2_11),
                        .Slide_data_12(in_data_to_next_pe_2_12), .Slide_data_13(in_data_to_next_pe_2_13),
                        .Slide_data_14(in_data_to_next_pe_2_14), .Slide_data_15(in_data_to_next_pe_2_15),
                        .Slide_data_16(in_data_to_next_pe_2_16), .Slide_data_17(in_data_to_next_pe_2_17),
                        .Slide_data_18(in_data_to_next_pe_2_18), .Slide_data_19(in_data_to_next_pe_2_19),
                        .Slide_data_20(in_data_to_next_pe_2_20), .Slide_data_21(in_data_to_next_pe_2_21),
                        .Slide_data_22(in_data_to_next_pe_2_22), .Slide_data_23(in_data_to_next_pe_2_23),
                        .Slide_data_24(in_data_to_next_pe_2_24), .Slide_data_25(in_data_to_next_pe_2_25),
                        .Slide_data_26(in_data_to_next_pe_2_26), .Slide_data_27(in_data_to_next_pe_2_27),
                        .Slide_data_28(in_data_to_next_pe_2_28), .Slide_data_29(in_data_to_next_pe_2_29),
                        .Slide_data_30(in_data_to_next_pe_2_30), .Slide_data_31(in_data_to_next_pe_2_31),
                        .result(o_2),
                        .in_data_to_next_pe_0(in_data_to_next_pe_3_0), .in_data_to_next_pe_1(in_data_to_next_pe_3_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_3_2), .in_data_to_next_pe_3(in_data_to_next_pe_3_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_3_4), .in_data_to_next_pe_5(in_data_to_next_pe_3_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_3_6), .in_data_to_next_pe_7(in_data_to_next_pe_3_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_3_8), .in_data_to_next_pe_9(in_data_to_next_pe_3_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_3_10), .in_data_to_next_pe_11(in_data_to_next_pe_3_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_3_12), .in_data_to_next_pe_13(in_data_to_next_pe_3_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_3_14), .in_data_to_next_pe_15(in_data_to_next_pe_3_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_3_16), .in_data_to_next_pe_17(in_data_to_next_pe_3_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_3_18), .in_data_to_next_pe_19(in_data_to_next_pe_3_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_3_20), .in_data_to_next_pe_21(in_data_to_next_pe_3_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_3_22), .in_data_to_next_pe_23(in_data_to_next_pe_3_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_3_24), .in_data_to_next_pe_25(in_data_to_next_pe_3_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_3_26), .in_data_to_next_pe_27(in_data_to_next_pe_3_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_3_28), .in_data_to_next_pe_29(in_data_to_next_pe_3_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_3_30), .in_data_to_next_pe_31(in_data_to_next_pe_3_31),
                        .next_row_en(row_3_en)
        );
        
        PE_Row_B5   PE_R3_B5(   .clk(clk), .rst_n(row_3_en), .new_weight_val(new_weight_val[3]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_3_0), .Slide_data_1(in_data_to_next_pe_3_1),
                        .Slide_data_2(in_data_to_next_pe_3_2), .Slide_data_3(in_data_to_next_pe_3_3),
                        .Slide_data_4(in_data_to_next_pe_3_4), .Slide_data_5(in_data_to_next_pe_3_5),
                        .Slide_data_6(in_data_to_next_pe_3_6), .Slide_data_7(in_data_to_next_pe_3_7),
                        .Slide_data_8(in_data_to_next_pe_3_8), .Slide_data_9(in_data_to_next_pe_3_9),
                        .Slide_data_10(in_data_to_next_pe_3_10), .Slide_data_11(in_data_to_next_pe_3_11),
                        .Slide_data_12(in_data_to_next_pe_3_12), .Slide_data_13(in_data_to_next_pe_3_13),
                        .Slide_data_14(in_data_to_next_pe_3_14), .Slide_data_15(in_data_to_next_pe_3_15),
                        .Slide_data_16(in_data_to_next_pe_3_16), .Slide_data_17(in_data_to_next_pe_3_17),
                        .Slide_data_18(in_data_to_next_pe_3_18), .Slide_data_19(in_data_to_next_pe_3_19),
                        .Slide_data_20(in_data_to_next_pe_3_20), .Slide_data_21(in_data_to_next_pe_3_21),
                        .Slide_data_22(in_data_to_next_pe_3_22), .Slide_data_23(in_data_to_next_pe_3_23),
                        .Slide_data_24(in_data_to_next_pe_3_24), .Slide_data_25(in_data_to_next_pe_3_25),
                        .Slide_data_26(in_data_to_next_pe_3_26), .Slide_data_27(in_data_to_next_pe_3_27),
                        .Slide_data_28(in_data_to_next_pe_3_28), .Slide_data_29(in_data_to_next_pe_3_29),
                        .Slide_data_30(in_data_to_next_pe_3_30), .Slide_data_31(in_data_to_next_pe_3_31),
                        .result(o_3),
                        .in_data_to_next_pe_0(in_data_to_next_pe_4_0), .in_data_to_next_pe_1(in_data_to_next_pe_4_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_4_2), .in_data_to_next_pe_3(in_data_to_next_pe_4_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_4_4), .in_data_to_next_pe_5(in_data_to_next_pe_4_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_4_6), .in_data_to_next_pe_7(in_data_to_next_pe_4_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_4_8), .in_data_to_next_pe_9(in_data_to_next_pe_4_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_4_10), .in_data_to_next_pe_11(in_data_to_next_pe_4_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_4_12), .in_data_to_next_pe_13(in_data_to_next_pe_4_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_4_14), .in_data_to_next_pe_15(in_data_to_next_pe_4_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_4_16), .in_data_to_next_pe_17(in_data_to_next_pe_4_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_4_18), .in_data_to_next_pe_19(in_data_to_next_pe_4_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_4_20), .in_data_to_next_pe_21(in_data_to_next_pe_4_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_4_22), .in_data_to_next_pe_23(in_data_to_next_pe_4_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_4_24), .in_data_to_next_pe_25(in_data_to_next_pe_4_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_4_26), .in_data_to_next_pe_27(in_data_to_next_pe_4_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_4_28), .in_data_to_next_pe_29(in_data_to_next_pe_4_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_4_30), .in_data_to_next_pe_31(in_data_to_next_pe_4_31),
                        .next_row_en(row_4_en)
        );
        
        PE_Row_B5   PE_R4_B5(   .clk(clk), .rst_n(row_4_en), .new_weight_val(new_weight_val[4]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_4_0), .Slide_data_1(in_data_to_next_pe_4_1),
                        .Slide_data_2(in_data_to_next_pe_4_2), .Slide_data_3(in_data_to_next_pe_4_3),
                        .Slide_data_4(in_data_to_next_pe_4_4), .Slide_data_5(in_data_to_next_pe_4_5),
                        .Slide_data_6(in_data_to_next_pe_4_6), .Slide_data_7(in_data_to_next_pe_4_7),
                        .Slide_data_8(in_data_to_next_pe_4_8), .Slide_data_9(in_data_to_next_pe_4_9),
                        .Slide_data_10(in_data_to_next_pe_4_10), .Slide_data_11(in_data_to_next_pe_4_11),
                        .Slide_data_12(in_data_to_next_pe_4_12), .Slide_data_13(in_data_to_next_pe_4_13),
                        .Slide_data_14(in_data_to_next_pe_4_14), .Slide_data_15(in_data_to_next_pe_4_15),
                        .Slide_data_16(in_data_to_next_pe_4_16), .Slide_data_17(in_data_to_next_pe_4_17),
                        .Slide_data_18(in_data_to_next_pe_4_18), .Slide_data_19(in_data_to_next_pe_4_19),
                        .Slide_data_20(in_data_to_next_pe_4_20), .Slide_data_21(in_data_to_next_pe_4_21),
                        .Slide_data_22(in_data_to_next_pe_4_22), .Slide_data_23(in_data_to_next_pe_4_23),
                        .Slide_data_24(in_data_to_next_pe_4_24), .Slide_data_25(in_data_to_next_pe_4_25),
                        .Slide_data_26(in_data_to_next_pe_4_26), .Slide_data_27(in_data_to_next_pe_4_27),
                        .Slide_data_28(in_data_to_next_pe_4_28), .Slide_data_29(in_data_to_next_pe_4_29),
                        .Slide_data_30(in_data_to_next_pe_4_30), .Slide_data_31(in_data_to_next_pe_4_31),
                        .result(o_4),
                        .in_data_to_next_pe_0(in_data_to_next_pe_5_0), .in_data_to_next_pe_1(in_data_to_next_pe_5_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_5_2), .in_data_to_next_pe_3(in_data_to_next_pe_5_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_5_4), .in_data_to_next_pe_5(in_data_to_next_pe_5_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_5_6), .in_data_to_next_pe_7(in_data_to_next_pe_5_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_5_8), .in_data_to_next_pe_9(in_data_to_next_pe_5_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_5_10), .in_data_to_next_pe_11(in_data_to_next_pe_5_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_5_12), .in_data_to_next_pe_13(in_data_to_next_pe_5_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_5_14), .in_data_to_next_pe_15(in_data_to_next_pe_5_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_5_16), .in_data_to_next_pe_17(in_data_to_next_pe_5_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_5_18), .in_data_to_next_pe_19(in_data_to_next_pe_5_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_5_20), .in_data_to_next_pe_21(in_data_to_next_pe_5_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_5_22), .in_data_to_next_pe_23(in_data_to_next_pe_5_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_5_24), .in_data_to_next_pe_25(in_data_to_next_pe_5_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_5_26), .in_data_to_next_pe_27(in_data_to_next_pe_5_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_5_28), .in_data_to_next_pe_29(in_data_to_next_pe_5_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_5_30), .in_data_to_next_pe_31(in_data_to_next_pe_5_31),
                        .next_row_en(row_5_en)
        );
        
        PE_Row_B5   PE_R5_B5(   .clk(clk), .rst_n(row_5_en), .new_weight_val(new_weight_val[5]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_5_0), .Slide_data_1(in_data_to_next_pe_5_1),
                        .Slide_data_2(in_data_to_next_pe_5_2), .Slide_data_3(in_data_to_next_pe_5_3),
                        .Slide_data_4(in_data_to_next_pe_5_4), .Slide_data_5(in_data_to_next_pe_5_5),
                        .Slide_data_6(in_data_to_next_pe_5_6), .Slide_data_7(in_data_to_next_pe_5_7),
                        .Slide_data_8(in_data_to_next_pe_5_8), .Slide_data_9(in_data_to_next_pe_5_9),
                        .Slide_data_10(in_data_to_next_pe_5_10), .Slide_data_11(in_data_to_next_pe_5_11),
                        .Slide_data_12(in_data_to_next_pe_5_12), .Slide_data_13(in_data_to_next_pe_5_13),
                        .Slide_data_14(in_data_to_next_pe_5_14), .Slide_data_15(in_data_to_next_pe_5_15),
                        .Slide_data_16(in_data_to_next_pe_5_16), .Slide_data_17(in_data_to_next_pe_5_17),
                        .Slide_data_18(in_data_to_next_pe_5_18), .Slide_data_19(in_data_to_next_pe_5_19),
                        .Slide_data_20(in_data_to_next_pe_5_20), .Slide_data_21(in_data_to_next_pe_5_21),
                        .Slide_data_22(in_data_to_next_pe_5_22), .Slide_data_23(in_data_to_next_pe_5_23),
                        .Slide_data_24(in_data_to_next_pe_5_24), .Slide_data_25(in_data_to_next_pe_5_25),
                        .Slide_data_26(in_data_to_next_pe_5_26), .Slide_data_27(in_data_to_next_pe_5_27),
                        .Slide_data_28(in_data_to_next_pe_5_28), .Slide_data_29(in_data_to_next_pe_5_29),
                        .Slide_data_30(in_data_to_next_pe_5_30), .Slide_data_31(in_data_to_next_pe_5_31),
                        .result(o_5),
                        .in_data_to_next_pe_0(in_data_to_next_pe_6_0), .in_data_to_next_pe_1(in_data_to_next_pe_6_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_6_2), .in_data_to_next_pe_3(in_data_to_next_pe_6_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_6_4), .in_data_to_next_pe_5(in_data_to_next_pe_6_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_6_6), .in_data_to_next_pe_7(in_data_to_next_pe_6_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_6_8), .in_data_to_next_pe_9(in_data_to_next_pe_6_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_6_10), .in_data_to_next_pe_11(in_data_to_next_pe_6_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_6_12), .in_data_to_next_pe_13(in_data_to_next_pe_6_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_6_14), .in_data_to_next_pe_15(in_data_to_next_pe_6_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_6_16), .in_data_to_next_pe_17(in_data_to_next_pe_6_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_6_18), .in_data_to_next_pe_19(in_data_to_next_pe_6_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_6_20), .in_data_to_next_pe_21(in_data_to_next_pe_6_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_6_22), .in_data_to_next_pe_23(in_data_to_next_pe_6_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_6_24), .in_data_to_next_pe_25(in_data_to_next_pe_6_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_6_26), .in_data_to_next_pe_27(in_data_to_next_pe_6_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_6_28), .in_data_to_next_pe_29(in_data_to_next_pe_6_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_6_30), .in_data_to_next_pe_31(in_data_to_next_pe_6_31),
                        .next_row_en(row_6_en)
        );
        
        PE_Row_B5   PE_R6_B5(   .clk(clk), .rst_n(row_6_en), .new_weight_val(new_weight_val[6]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_6_0), .Slide_data_1(in_data_to_next_pe_6_1),
                        .Slide_data_2(in_data_to_next_pe_6_2), .Slide_data_3(in_data_to_next_pe_6_3),
                        .Slide_data_4(in_data_to_next_pe_6_4), .Slide_data_5(in_data_to_next_pe_6_5),
                        .Slide_data_6(in_data_to_next_pe_6_6), .Slide_data_7(in_data_to_next_pe_6_7),
                        .Slide_data_8(in_data_to_next_pe_6_8), .Slide_data_9(in_data_to_next_pe_6_9),
                        .Slide_data_10(in_data_to_next_pe_6_10), .Slide_data_11(in_data_to_next_pe_6_11),
                        .Slide_data_12(in_data_to_next_pe_6_12), .Slide_data_13(in_data_to_next_pe_6_13),
                        .Slide_data_14(in_data_to_next_pe_6_14), .Slide_data_15(in_data_to_next_pe_6_15),
                        .Slide_data_16(in_data_to_next_pe_6_16), .Slide_data_17(in_data_to_next_pe_6_17),
                        .Slide_data_18(in_data_to_next_pe_6_18), .Slide_data_19(in_data_to_next_pe_6_19),
                        .Slide_data_20(in_data_to_next_pe_6_20), .Slide_data_21(in_data_to_next_pe_6_21),
                        .Slide_data_22(in_data_to_next_pe_6_22), .Slide_data_23(in_data_to_next_pe_6_23),
                        .Slide_data_24(in_data_to_next_pe_6_24), .Slide_data_25(in_data_to_next_pe_6_25),
                        .Slide_data_26(in_data_to_next_pe_6_26), .Slide_data_27(in_data_to_next_pe_6_27),
                        .Slide_data_28(in_data_to_next_pe_6_28), .Slide_data_29(in_data_to_next_pe_6_29),
                        .Slide_data_30(in_data_to_next_pe_6_30), .Slide_data_31(in_data_to_next_pe_6_31),
                        .result(o_6),
                        .in_data_to_next_pe_0(in_data_to_next_pe_7_0), .in_data_to_next_pe_1(in_data_to_next_pe_7_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_7_2), .in_data_to_next_pe_3(in_data_to_next_pe_7_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_7_4), .in_data_to_next_pe_5(in_data_to_next_pe_7_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_7_6), .in_data_to_next_pe_7(in_data_to_next_pe_7_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_7_8), .in_data_to_next_pe_9(in_data_to_next_pe_7_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_7_10), .in_data_to_next_pe_11(in_data_to_next_pe_7_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_7_12), .in_data_to_next_pe_13(in_data_to_next_pe_7_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_7_14), .in_data_to_next_pe_15(in_data_to_next_pe_7_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_7_16), .in_data_to_next_pe_17(in_data_to_next_pe_7_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_7_18), .in_data_to_next_pe_19(in_data_to_next_pe_7_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_7_20), .in_data_to_next_pe_21(in_data_to_next_pe_7_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_7_22), .in_data_to_next_pe_23(in_data_to_next_pe_7_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_7_24), .in_data_to_next_pe_25(in_data_to_next_pe_7_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_7_26), .in_data_to_next_pe_27(in_data_to_next_pe_7_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_7_28), .in_data_to_next_pe_29(in_data_to_next_pe_7_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_7_30), .in_data_to_next_pe_31(in_data_to_next_pe_7_31),
                        .next_row_en(row_7_en)
        );
        
        PE_Row_B5   PE_R7_B5(   .clk(clk), .rst_n(row_7_en), .new_weight_val(new_weight_val[7]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_7_0), .Slide_data_1(in_data_to_next_pe_7_1),
                        .Slide_data_2(in_data_to_next_pe_7_2), .Slide_data_3(in_data_to_next_pe_7_3),
                        .Slide_data_4(in_data_to_next_pe_7_4), .Slide_data_5(in_data_to_next_pe_7_5),
                        .Slide_data_6(in_data_to_next_pe_7_6), .Slide_data_7(in_data_to_next_pe_7_7),
                        .Slide_data_8(in_data_to_next_pe_7_8), .Slide_data_9(in_data_to_next_pe_7_9),
                        .Slide_data_10(in_data_to_next_pe_7_10), .Slide_data_11(in_data_to_next_pe_7_11),
                        .Slide_data_12(in_data_to_next_pe_7_12), .Slide_data_13(in_data_to_next_pe_7_13),
                        .Slide_data_14(in_data_to_next_pe_7_14), .Slide_data_15(in_data_to_next_pe_7_15),
                        .Slide_data_16(in_data_to_next_pe_7_16), .Slide_data_17(in_data_to_next_pe_7_17),
                        .Slide_data_18(in_data_to_next_pe_7_18), .Slide_data_19(in_data_to_next_pe_7_19),
                        .Slide_data_20(in_data_to_next_pe_7_20), .Slide_data_21(in_data_to_next_pe_7_21),
                        .Slide_data_22(in_data_to_next_pe_7_22), .Slide_data_23(in_data_to_next_pe_7_23),
                        .Slide_data_24(in_data_to_next_pe_7_24), .Slide_data_25(in_data_to_next_pe_7_25),
                        .Slide_data_26(in_data_to_next_pe_7_26), .Slide_data_27(in_data_to_next_pe_7_27),
                        .Slide_data_28(in_data_to_next_pe_7_28), .Slide_data_29(in_data_to_next_pe_7_29),
                        .Slide_data_30(in_data_to_next_pe_7_30), .Slide_data_31(in_data_to_next_pe_7_31),
                        .result(o_7),
                        .in_data_to_next_pe_0(in_data_to_next_pe_8_0), .in_data_to_next_pe_1(in_data_to_next_pe_8_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_8_2), .in_data_to_next_pe_3(in_data_to_next_pe_8_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_8_4), .in_data_to_next_pe_5(in_data_to_next_pe_8_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_8_6), .in_data_to_next_pe_7(in_data_to_next_pe_8_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_8_8), .in_data_to_next_pe_9(in_data_to_next_pe_8_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_8_10), .in_data_to_next_pe_11(in_data_to_next_pe_8_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_8_12), .in_data_to_next_pe_13(in_data_to_next_pe_8_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_8_14), .in_data_to_next_pe_15(in_data_to_next_pe_8_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_8_16), .in_data_to_next_pe_17(in_data_to_next_pe_8_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_8_18), .in_data_to_next_pe_19(in_data_to_next_pe_8_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_8_20), .in_data_to_next_pe_21(in_data_to_next_pe_8_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_8_22), .in_data_to_next_pe_23(in_data_to_next_pe_8_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_8_24), .in_data_to_next_pe_25(in_data_to_next_pe_8_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_8_26), .in_data_to_next_pe_27(in_data_to_next_pe_8_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_8_28), .in_data_to_next_pe_29(in_data_to_next_pe_8_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_8_30), .in_data_to_next_pe_31(in_data_to_next_pe_8_31),
                        .next_row_en(row_8_en)
        );
        
        PE_Row_B5   PE_R8_B5(   .clk(clk), .rst_n(row_8_en), .new_weight_val(new_weight_val[8]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_8_0), .Slide_data_1(in_data_to_next_pe_8_1),
                        .Slide_data_2(in_data_to_next_pe_8_2), .Slide_data_3(in_data_to_next_pe_8_3),
                        .Slide_data_4(in_data_to_next_pe_8_4), .Slide_data_5(in_data_to_next_pe_8_5),
                        .Slide_data_6(in_data_to_next_pe_8_6), .Slide_data_7(in_data_to_next_pe_8_7),
                        .Slide_data_8(in_data_to_next_pe_8_8), .Slide_data_9(in_data_to_next_pe_8_9),
                        .Slide_data_10(in_data_to_next_pe_8_10), .Slide_data_11(in_data_to_next_pe_8_11),
                        .Slide_data_12(in_data_to_next_pe_8_12), .Slide_data_13(in_data_to_next_pe_8_13),
                        .Slide_data_14(in_data_to_next_pe_8_14), .Slide_data_15(in_data_to_next_pe_8_15),
                        .Slide_data_16(in_data_to_next_pe_8_16), .Slide_data_17(in_data_to_next_pe_8_17),
                        .Slide_data_18(in_data_to_next_pe_8_18), .Slide_data_19(in_data_to_next_pe_8_19),
                        .Slide_data_20(in_data_to_next_pe_8_20), .Slide_data_21(in_data_to_next_pe_8_21),
                        .Slide_data_22(in_data_to_next_pe_8_22), .Slide_data_23(in_data_to_next_pe_8_23),
                        .Slide_data_24(in_data_to_next_pe_8_24), .Slide_data_25(in_data_to_next_pe_8_25),
                        .Slide_data_26(in_data_to_next_pe_8_26), .Slide_data_27(in_data_to_next_pe_8_27),
                        .Slide_data_28(in_data_to_next_pe_8_28), .Slide_data_29(in_data_to_next_pe_8_29),
                        .Slide_data_30(in_data_to_next_pe_8_30), .Slide_data_31(in_data_to_next_pe_8_31),
                        .result(o_8),
                        .in_data_to_next_pe_0(in_data_to_next_pe_9_0), .in_data_to_next_pe_1(in_data_to_next_pe_9_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_9_2), .in_data_to_next_pe_3(in_data_to_next_pe_9_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_9_4), .in_data_to_next_pe_5(in_data_to_next_pe_9_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_9_6), .in_data_to_next_pe_7(in_data_to_next_pe_9_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_9_8), .in_data_to_next_pe_9(in_data_to_next_pe_9_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_9_10), .in_data_to_next_pe_11(in_data_to_next_pe_9_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_9_12), .in_data_to_next_pe_13(in_data_to_next_pe_9_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_9_14), .in_data_to_next_pe_15(in_data_to_next_pe_9_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_9_16), .in_data_to_next_pe_17(in_data_to_next_pe_9_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_9_18), .in_data_to_next_pe_19(in_data_to_next_pe_9_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_9_20), .in_data_to_next_pe_21(in_data_to_next_pe_9_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_9_22), .in_data_to_next_pe_23(in_data_to_next_pe_9_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_9_24), .in_data_to_next_pe_25(in_data_to_next_pe_9_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_9_26), .in_data_to_next_pe_27(in_data_to_next_pe_9_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_9_28), .in_data_to_next_pe_29(in_data_to_next_pe_9_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_9_30), .in_data_to_next_pe_31(in_data_to_next_pe_9_31),
                        .next_row_en(row_9_en)
        );
        
        PE_Row_B5   PE_R9_B5(   .clk(clk), .rst_n(row_9_en), .new_weight_val(new_weight_val[9]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_9_0), .Slide_data_1(in_data_to_next_pe_9_1),
                        .Slide_data_2(in_data_to_next_pe_9_2), .Slide_data_3(in_data_to_next_pe_9_3),
                        .Slide_data_4(in_data_to_next_pe_9_4), .Slide_data_5(in_data_to_next_pe_9_5),
                        .Slide_data_6(in_data_to_next_pe_9_6), .Slide_data_7(in_data_to_next_pe_9_7),
                        .Slide_data_8(in_data_to_next_pe_9_8), .Slide_data_9(in_data_to_next_pe_9_9),
                        .Slide_data_10(in_data_to_next_pe_9_10), .Slide_data_11(in_data_to_next_pe_9_11),
                        .Slide_data_12(in_data_to_next_pe_9_12), .Slide_data_13(in_data_to_next_pe_9_13),
                        .Slide_data_14(in_data_to_next_pe_9_14), .Slide_data_15(in_data_to_next_pe_9_15),
                        .Slide_data_16(in_data_to_next_pe_9_16), .Slide_data_17(in_data_to_next_pe_9_17),
                        .Slide_data_18(in_data_to_next_pe_9_18), .Slide_data_19(in_data_to_next_pe_9_19),
                        .Slide_data_20(in_data_to_next_pe_9_20), .Slide_data_21(in_data_to_next_pe_9_21),
                        .Slide_data_22(in_data_to_next_pe_9_22), .Slide_data_23(in_data_to_next_pe_9_23),
                        .Slide_data_24(in_data_to_next_pe_9_24), .Slide_data_25(in_data_to_next_pe_9_25),
                        .Slide_data_26(in_data_to_next_pe_9_26), .Slide_data_27(in_data_to_next_pe_9_27),
                        .Slide_data_28(in_data_to_next_pe_9_28), .Slide_data_29(in_data_to_next_pe_9_29),
                        .Slide_data_30(in_data_to_next_pe_9_30), .Slide_data_31(in_data_to_next_pe_9_31),
                        .result(o_9),
                        .in_data_to_next_pe_0(in_data_to_next_pe_10_0), .in_data_to_next_pe_1(in_data_to_next_pe_10_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_10_2), .in_data_to_next_pe_3(in_data_to_next_pe_10_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_10_4), .in_data_to_next_pe_5(in_data_to_next_pe_10_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_10_6), .in_data_to_next_pe_7(in_data_to_next_pe_10_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_10_8), .in_data_to_next_pe_9(in_data_to_next_pe_10_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_10_10), .in_data_to_next_pe_11(in_data_to_next_pe_10_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_10_12), .in_data_to_next_pe_13(in_data_to_next_pe_10_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_10_14), .in_data_to_next_pe_15(in_data_to_next_pe_10_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_10_16), .in_data_to_next_pe_17(in_data_to_next_pe_10_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_10_18), .in_data_to_next_pe_19(in_data_to_next_pe_10_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_10_20), .in_data_to_next_pe_21(in_data_to_next_pe_10_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_10_22), .in_data_to_next_pe_23(in_data_to_next_pe_10_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_10_24), .in_data_to_next_pe_25(in_data_to_next_pe_10_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_10_26), .in_data_to_next_pe_27(in_data_to_next_pe_10_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_10_28), .in_data_to_next_pe_29(in_data_to_next_pe_10_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_10_30), .in_data_to_next_pe_31(in_data_to_next_pe_10_31),
                        .next_row_en(row_10_en)
        );
        
        PE_Row_B5   PE_R10_B5(   .clk(clk), .rst_n(row_10_en), .new_weight_val(new_weight_val[10]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_10_0), .Slide_data_1(in_data_to_next_pe_10_1),
                        .Slide_data_2(in_data_to_next_pe_10_2), .Slide_data_3(in_data_to_next_pe_10_3),
                        .Slide_data_4(in_data_to_next_pe_10_4), .Slide_data_5(in_data_to_next_pe_10_5),
                        .Slide_data_6(in_data_to_next_pe_10_6), .Slide_data_7(in_data_to_next_pe_10_7),
                        .Slide_data_8(in_data_to_next_pe_10_8), .Slide_data_9(in_data_to_next_pe_10_9),
                        .Slide_data_10(in_data_to_next_pe_10_10), .Slide_data_11(in_data_to_next_pe_10_11),
                        .Slide_data_12(in_data_to_next_pe_10_12), .Slide_data_13(in_data_to_next_pe_10_13),
                        .Slide_data_14(in_data_to_next_pe_10_14), .Slide_data_15(in_data_to_next_pe_10_15),
                        .Slide_data_16(in_data_to_next_pe_10_16), .Slide_data_17(in_data_to_next_pe_10_17),
                        .Slide_data_18(in_data_to_next_pe_10_18), .Slide_data_19(in_data_to_next_pe_10_19),
                        .Slide_data_20(in_data_to_next_pe_10_20), .Slide_data_21(in_data_to_next_pe_10_21),
                        .Slide_data_22(in_data_to_next_pe_10_22), .Slide_data_23(in_data_to_next_pe_10_23),
                        .Slide_data_24(in_data_to_next_pe_10_24), .Slide_data_25(in_data_to_next_pe_10_25),
                        .Slide_data_26(in_data_to_next_pe_10_26), .Slide_data_27(in_data_to_next_pe_10_27),
                        .Slide_data_28(in_data_to_next_pe_10_28), .Slide_data_29(in_data_to_next_pe_10_29),
                        .Slide_data_30(in_data_to_next_pe_10_30), .Slide_data_31(in_data_to_next_pe_10_31),
                        .result(o_10),
                        .in_data_to_next_pe_0(in_data_to_next_pe_11_0), .in_data_to_next_pe_1(in_data_to_next_pe_11_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_11_2), .in_data_to_next_pe_3(in_data_to_next_pe_11_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_11_4), .in_data_to_next_pe_5(in_data_to_next_pe_11_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_11_6), .in_data_to_next_pe_7(in_data_to_next_pe_11_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_11_8), .in_data_to_next_pe_9(in_data_to_next_pe_11_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_11_10), .in_data_to_next_pe_11(in_data_to_next_pe_11_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_11_12), .in_data_to_next_pe_13(in_data_to_next_pe_11_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_11_14), .in_data_to_next_pe_15(in_data_to_next_pe_11_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_11_16), .in_data_to_next_pe_17(in_data_to_next_pe_11_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_11_18), .in_data_to_next_pe_19(in_data_to_next_pe_11_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_11_20), .in_data_to_next_pe_21(in_data_to_next_pe_11_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_11_22), .in_data_to_next_pe_23(in_data_to_next_pe_11_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_11_24), .in_data_to_next_pe_25(in_data_to_next_pe_11_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_11_26), .in_data_to_next_pe_27(in_data_to_next_pe_11_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_11_28), .in_data_to_next_pe_29(in_data_to_next_pe_11_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_11_30), .in_data_to_next_pe_31(in_data_to_next_pe_11_31),
                        .next_row_en(row_11_en)
        );
        
        PE_Row_B5   PE_R11_B5(   .clk(clk), .rst_n(row_11_en), .new_weight_val(new_weight_val[11]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_11_0), .Slide_data_1(in_data_to_next_pe_11_1),
                        .Slide_data_2(in_data_to_next_pe_11_2), .Slide_data_3(in_data_to_next_pe_11_3),
                        .Slide_data_4(in_data_to_next_pe_11_4), .Slide_data_5(in_data_to_next_pe_11_5),
                        .Slide_data_6(in_data_to_next_pe_11_6), .Slide_data_7(in_data_to_next_pe_11_7),
                        .Slide_data_8(in_data_to_next_pe_11_8), .Slide_data_9(in_data_to_next_pe_11_9),
                        .Slide_data_10(in_data_to_next_pe_11_10), .Slide_data_11(in_data_to_next_pe_11_11),
                        .Slide_data_12(in_data_to_next_pe_11_12), .Slide_data_13(in_data_to_next_pe_11_13),
                        .Slide_data_14(in_data_to_next_pe_11_14), .Slide_data_15(in_data_to_next_pe_11_15),
                        .Slide_data_16(in_data_to_next_pe_11_16), .Slide_data_17(in_data_to_next_pe_11_17),
                        .Slide_data_18(in_data_to_next_pe_11_18), .Slide_data_19(in_data_to_next_pe_11_19),
                        .Slide_data_20(in_data_to_next_pe_11_20), .Slide_data_21(in_data_to_next_pe_11_21),
                        .Slide_data_22(in_data_to_next_pe_11_22), .Slide_data_23(in_data_to_next_pe_11_23),
                        .Slide_data_24(in_data_to_next_pe_11_24), .Slide_data_25(in_data_to_next_pe_11_25),
                        .Slide_data_26(in_data_to_next_pe_11_26), .Slide_data_27(in_data_to_next_pe_11_27),
                        .Slide_data_28(in_data_to_next_pe_11_28), .Slide_data_29(in_data_to_next_pe_11_29),
                        .Slide_data_30(in_data_to_next_pe_11_30), .Slide_data_31(in_data_to_next_pe_11_31),
                        .result(o_11),
                        .in_data_to_next_pe_0(in_data_to_next_pe_12_0), .in_data_to_next_pe_1(in_data_to_next_pe_12_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_12_2), .in_data_to_next_pe_3(in_data_to_next_pe_12_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_12_4), .in_data_to_next_pe_5(in_data_to_next_pe_12_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_12_6), .in_data_to_next_pe_7(in_data_to_next_pe_12_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_12_8), .in_data_to_next_pe_9(in_data_to_next_pe_12_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_12_10), .in_data_to_next_pe_11(in_data_to_next_pe_12_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_12_12), .in_data_to_next_pe_13(in_data_to_next_pe_12_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_12_14), .in_data_to_next_pe_15(in_data_to_next_pe_12_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_12_16), .in_data_to_next_pe_17(in_data_to_next_pe_12_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_12_18), .in_data_to_next_pe_19(in_data_to_next_pe_12_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_12_20), .in_data_to_next_pe_21(in_data_to_next_pe_12_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_12_22), .in_data_to_next_pe_23(in_data_to_next_pe_12_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_12_24), .in_data_to_next_pe_25(in_data_to_next_pe_12_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_12_26), .in_data_to_next_pe_27(in_data_to_next_pe_12_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_12_28), .in_data_to_next_pe_29(in_data_to_next_pe_12_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_12_30), .in_data_to_next_pe_31(in_data_to_next_pe_12_31),
                        .next_row_en(row_12_en)
        );
        
        PE_Row_B5   PE_R12_B5(   .clk(clk), .rst_n(row_12_en), .new_weight_val(new_weight_val[12]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_12_0), .Slide_data_1(in_data_to_next_pe_12_1),
                        .Slide_data_2(in_data_to_next_pe_12_2), .Slide_data_3(in_data_to_next_pe_12_3),
                        .Slide_data_4(in_data_to_next_pe_12_4), .Slide_data_5(in_data_to_next_pe_12_5),
                        .Slide_data_6(in_data_to_next_pe_12_6), .Slide_data_7(in_data_to_next_pe_12_7),
                        .Slide_data_8(in_data_to_next_pe_12_8), .Slide_data_9(in_data_to_next_pe_12_9),
                        .Slide_data_10(in_data_to_next_pe_12_10), .Slide_data_11(in_data_to_next_pe_12_11),
                        .Slide_data_12(in_data_to_next_pe_12_12), .Slide_data_13(in_data_to_next_pe_12_13),
                        .Slide_data_14(in_data_to_next_pe_12_14), .Slide_data_15(in_data_to_next_pe_12_15),
                        .Slide_data_16(in_data_to_next_pe_12_16), .Slide_data_17(in_data_to_next_pe_12_17),
                        .Slide_data_18(in_data_to_next_pe_12_18), .Slide_data_19(in_data_to_next_pe_12_19),
                        .Slide_data_20(in_data_to_next_pe_12_20), .Slide_data_21(in_data_to_next_pe_12_21),
                        .Slide_data_22(in_data_to_next_pe_12_22), .Slide_data_23(in_data_to_next_pe_12_23),
                        .Slide_data_24(in_data_to_next_pe_12_24), .Slide_data_25(in_data_to_next_pe_12_25),
                        .Slide_data_26(in_data_to_next_pe_12_26), .Slide_data_27(in_data_to_next_pe_12_27),
                        .Slide_data_28(in_data_to_next_pe_12_28), .Slide_data_29(in_data_to_next_pe_12_29),
                        .Slide_data_30(in_data_to_next_pe_12_30), .Slide_data_31(in_data_to_next_pe_12_31),
                        .result(o_12),
                        .in_data_to_next_pe_0(in_data_to_next_pe_13_0), .in_data_to_next_pe_1(in_data_to_next_pe_13_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_13_2), .in_data_to_next_pe_3(in_data_to_next_pe_13_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_13_4), .in_data_to_next_pe_5(in_data_to_next_pe_13_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_13_6), .in_data_to_next_pe_7(in_data_to_next_pe_13_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_13_8), .in_data_to_next_pe_9(in_data_to_next_pe_13_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_13_10), .in_data_to_next_pe_11(in_data_to_next_pe_13_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_13_12), .in_data_to_next_pe_13(in_data_to_next_pe_13_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_13_14), .in_data_to_next_pe_15(in_data_to_next_pe_13_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_13_16), .in_data_to_next_pe_17(in_data_to_next_pe_13_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_13_18), .in_data_to_next_pe_19(in_data_to_next_pe_13_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_13_20), .in_data_to_next_pe_21(in_data_to_next_pe_13_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_13_22), .in_data_to_next_pe_23(in_data_to_next_pe_13_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_13_24), .in_data_to_next_pe_25(in_data_to_next_pe_13_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_13_26), .in_data_to_next_pe_27(in_data_to_next_pe_13_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_13_28), .in_data_to_next_pe_29(in_data_to_next_pe_13_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_13_30), .in_data_to_next_pe_31(in_data_to_next_pe_13_31),
                        .next_row_en(row_13_en)
        );
        
        PE_Row_B5   PE_R13_B5(   .clk(clk), .rst_n(row_13_en), .new_weight_val(new_weight_val[13]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_13_0), .Slide_data_1(in_data_to_next_pe_13_1),
                        .Slide_data_2(in_data_to_next_pe_13_2), .Slide_data_3(in_data_to_next_pe_13_3),
                        .Slide_data_4(in_data_to_next_pe_13_4), .Slide_data_5(in_data_to_next_pe_13_5),
                        .Slide_data_6(in_data_to_next_pe_13_6), .Slide_data_7(in_data_to_next_pe_13_7),
                        .Slide_data_8(in_data_to_next_pe_13_8), .Slide_data_9(in_data_to_next_pe_13_9),
                        .Slide_data_10(in_data_to_next_pe_13_10), .Slide_data_11(in_data_to_next_pe_13_11),
                        .Slide_data_12(in_data_to_next_pe_13_12), .Slide_data_13(in_data_to_next_pe_13_13),
                        .Slide_data_14(in_data_to_next_pe_13_14), .Slide_data_15(in_data_to_next_pe_13_15),
                        .Slide_data_16(in_data_to_next_pe_13_16), .Slide_data_17(in_data_to_next_pe_13_17),
                        .Slide_data_18(in_data_to_next_pe_13_18), .Slide_data_19(in_data_to_next_pe_13_19),
                        .Slide_data_20(in_data_to_next_pe_13_20), .Slide_data_21(in_data_to_next_pe_13_21),
                        .Slide_data_22(in_data_to_next_pe_13_22), .Slide_data_23(in_data_to_next_pe_13_23),
                        .Slide_data_24(in_data_to_next_pe_13_24), .Slide_data_25(in_data_to_next_pe_13_25),
                        .Slide_data_26(in_data_to_next_pe_13_26), .Slide_data_27(in_data_to_next_pe_13_27),
                        .Slide_data_28(in_data_to_next_pe_13_28), .Slide_data_29(in_data_to_next_pe_13_29),
                        .Slide_data_30(in_data_to_next_pe_13_30), .Slide_data_31(in_data_to_next_pe_13_31),
                        .result(o_13),
                        .in_data_to_next_pe_0(in_data_to_next_pe_14_0), .in_data_to_next_pe_1(in_data_to_next_pe_14_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_14_2), .in_data_to_next_pe_3(in_data_to_next_pe_14_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_14_4), .in_data_to_next_pe_5(in_data_to_next_pe_14_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_14_6), .in_data_to_next_pe_7(in_data_to_next_pe_14_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_14_8), .in_data_to_next_pe_9(in_data_to_next_pe_14_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_14_10), .in_data_to_next_pe_11(in_data_to_next_pe_14_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_14_12), .in_data_to_next_pe_13(in_data_to_next_pe_14_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_14_14), .in_data_to_next_pe_15(in_data_to_next_pe_14_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_14_16), .in_data_to_next_pe_17(in_data_to_next_pe_14_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_14_18), .in_data_to_next_pe_19(in_data_to_next_pe_14_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_14_20), .in_data_to_next_pe_21(in_data_to_next_pe_14_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_14_22), .in_data_to_next_pe_23(in_data_to_next_pe_14_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_14_24), .in_data_to_next_pe_25(in_data_to_next_pe_14_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_14_26), .in_data_to_next_pe_27(in_data_to_next_pe_14_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_14_28), .in_data_to_next_pe_29(in_data_to_next_pe_14_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_14_30), .in_data_to_next_pe_31(in_data_to_next_pe_14_31),
                        .next_row_en(row_14_en)
        );
        
        PE_Row_B5   PE_R14_B5(   .clk(clk), .rst_n(row_14_en), .new_weight_val(new_weight_val[14]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_14_0), .Slide_data_1(in_data_to_next_pe_14_1),
                        .Slide_data_2(in_data_to_next_pe_14_2), .Slide_data_3(in_data_to_next_pe_14_3),
                        .Slide_data_4(in_data_to_next_pe_14_4), .Slide_data_5(in_data_to_next_pe_14_5),
                        .Slide_data_6(in_data_to_next_pe_14_6), .Slide_data_7(in_data_to_next_pe_14_7),
                        .Slide_data_8(in_data_to_next_pe_14_8), .Slide_data_9(in_data_to_next_pe_14_9),
                        .Slide_data_10(in_data_to_next_pe_14_10), .Slide_data_11(in_data_to_next_pe_14_11),
                        .Slide_data_12(in_data_to_next_pe_14_12), .Slide_data_13(in_data_to_next_pe_14_13),
                        .Slide_data_14(in_data_to_next_pe_14_14), .Slide_data_15(in_data_to_next_pe_14_15),
                        .Slide_data_16(in_data_to_next_pe_14_16), .Slide_data_17(in_data_to_next_pe_14_17),
                        .Slide_data_18(in_data_to_next_pe_14_18), .Slide_data_19(in_data_to_next_pe_14_19),
                        .Slide_data_20(in_data_to_next_pe_14_20), .Slide_data_21(in_data_to_next_pe_14_21),
                        .Slide_data_22(in_data_to_next_pe_14_22), .Slide_data_23(in_data_to_next_pe_14_23),
                        .Slide_data_24(in_data_to_next_pe_14_24), .Slide_data_25(in_data_to_next_pe_14_25),
                        .Slide_data_26(in_data_to_next_pe_14_26), .Slide_data_27(in_data_to_next_pe_14_27),
                        .Slide_data_28(in_data_to_next_pe_14_28), .Slide_data_29(in_data_to_next_pe_14_29),
                        .Slide_data_30(in_data_to_next_pe_14_30), .Slide_data_31(in_data_to_next_pe_14_31),
                        .result(o_14),
                        .in_data_to_next_pe_0(in_data_to_next_pe_15_0), .in_data_to_next_pe_1(in_data_to_next_pe_15_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_15_2), .in_data_to_next_pe_3(in_data_to_next_pe_15_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_15_4), .in_data_to_next_pe_5(in_data_to_next_pe_15_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_15_6), .in_data_to_next_pe_7(in_data_to_next_pe_15_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_15_8), .in_data_to_next_pe_9(in_data_to_next_pe_15_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_15_10), .in_data_to_next_pe_11(in_data_to_next_pe_15_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_15_12), .in_data_to_next_pe_13(in_data_to_next_pe_15_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_15_14), .in_data_to_next_pe_15(in_data_to_next_pe_15_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_15_16), .in_data_to_next_pe_17(in_data_to_next_pe_15_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_15_18), .in_data_to_next_pe_19(in_data_to_next_pe_15_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_15_20), .in_data_to_next_pe_21(in_data_to_next_pe_15_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_15_22), .in_data_to_next_pe_23(in_data_to_next_pe_15_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_15_24), .in_data_to_next_pe_25(in_data_to_next_pe_15_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_15_26), .in_data_to_next_pe_27(in_data_to_next_pe_15_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_15_28), .in_data_to_next_pe_29(in_data_to_next_pe_15_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_15_30), .in_data_to_next_pe_31(in_data_to_next_pe_15_31),
                        .next_row_en(row_15_en)
        );
        
        PE_Row_B5   PE_R15_B5(   .clk(clk), .rst_n(row_15_en), .new_weight_val(new_weight_val[15]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_15_0), .Slide_data_1(in_data_to_next_pe_15_1),
                        .Slide_data_2(in_data_to_next_pe_15_2), .Slide_data_3(in_data_to_next_pe_15_3),
                        .Slide_data_4(in_data_to_next_pe_15_4), .Slide_data_5(in_data_to_next_pe_15_5),
                        .Slide_data_6(in_data_to_next_pe_15_6), .Slide_data_7(in_data_to_next_pe_15_7),
                        .Slide_data_8(in_data_to_next_pe_15_8), .Slide_data_9(in_data_to_next_pe_15_9),
                        .Slide_data_10(in_data_to_next_pe_15_10), .Slide_data_11(in_data_to_next_pe_15_11),
                        .Slide_data_12(in_data_to_next_pe_15_12), .Slide_data_13(in_data_to_next_pe_15_13),
                        .Slide_data_14(in_data_to_next_pe_15_14), .Slide_data_15(in_data_to_next_pe_15_15),
                        .Slide_data_16(in_data_to_next_pe_15_16), .Slide_data_17(in_data_to_next_pe_15_17),
                        .Slide_data_18(in_data_to_next_pe_15_18), .Slide_data_19(in_data_to_next_pe_15_19),
                        .Slide_data_20(in_data_to_next_pe_15_20), .Slide_data_21(in_data_to_next_pe_15_21),
                        .Slide_data_22(in_data_to_next_pe_15_22), .Slide_data_23(in_data_to_next_pe_15_23),
                        .Slide_data_24(in_data_to_next_pe_15_24), .Slide_data_25(in_data_to_next_pe_15_25),
                        .Slide_data_26(in_data_to_next_pe_15_26), .Slide_data_27(in_data_to_next_pe_15_27),
                        .Slide_data_28(in_data_to_next_pe_15_28), .Slide_data_29(in_data_to_next_pe_15_29),
                        .Slide_data_30(in_data_to_next_pe_15_30), .Slide_data_31(in_data_to_next_pe_15_31),
                        .result(o_15),
                        .in_data_to_next_pe_0(in_data_to_next_pe_16_0), .in_data_to_next_pe_1(in_data_to_next_pe_16_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_16_2), .in_data_to_next_pe_3(in_data_to_next_pe_16_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_16_4), .in_data_to_next_pe_5(in_data_to_next_pe_16_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_16_6), .in_data_to_next_pe_7(in_data_to_next_pe_16_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_16_8), .in_data_to_next_pe_9(in_data_to_next_pe_16_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_16_10), .in_data_to_next_pe_11(in_data_to_next_pe_16_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_16_12), .in_data_to_next_pe_13(in_data_to_next_pe_16_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_16_14), .in_data_to_next_pe_15(in_data_to_next_pe_16_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_16_16), .in_data_to_next_pe_17(in_data_to_next_pe_16_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_16_18), .in_data_to_next_pe_19(in_data_to_next_pe_16_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_16_20), .in_data_to_next_pe_21(in_data_to_next_pe_16_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_16_22), .in_data_to_next_pe_23(in_data_to_next_pe_16_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_16_24), .in_data_to_next_pe_25(in_data_to_next_pe_16_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_16_26), .in_data_to_next_pe_27(in_data_to_next_pe_16_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_16_28), .in_data_to_next_pe_29(in_data_to_next_pe_16_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_16_30), .in_data_to_next_pe_31(in_data_to_next_pe_16_31),
                        .next_row_en(row_16_en)
        );
        
        PE_Row_B5   PE_R16_B5(   .clk(clk), .rst_n(row_16_en), .new_weight_val(new_weight_val[16]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_16_0), .Slide_data_1(in_data_to_next_pe_16_1),
                        .Slide_data_2(in_data_to_next_pe_16_2), .Slide_data_3(in_data_to_next_pe_16_3),
                        .Slide_data_4(in_data_to_next_pe_16_4), .Slide_data_5(in_data_to_next_pe_16_5),
                        .Slide_data_6(in_data_to_next_pe_16_6), .Slide_data_7(in_data_to_next_pe_16_7),
                        .Slide_data_8(in_data_to_next_pe_16_8), .Slide_data_9(in_data_to_next_pe_16_9),
                        .Slide_data_10(in_data_to_next_pe_16_10), .Slide_data_11(in_data_to_next_pe_16_11),
                        .Slide_data_12(in_data_to_next_pe_16_12), .Slide_data_13(in_data_to_next_pe_16_13),
                        .Slide_data_14(in_data_to_next_pe_16_14), .Slide_data_15(in_data_to_next_pe_16_15),
                        .Slide_data_16(in_data_to_next_pe_16_16), .Slide_data_17(in_data_to_next_pe_16_17),
                        .Slide_data_18(in_data_to_next_pe_16_18), .Slide_data_19(in_data_to_next_pe_16_19),
                        .Slide_data_20(in_data_to_next_pe_16_20), .Slide_data_21(in_data_to_next_pe_16_21),
                        .Slide_data_22(in_data_to_next_pe_16_22), .Slide_data_23(in_data_to_next_pe_16_23),
                        .Slide_data_24(in_data_to_next_pe_16_24), .Slide_data_25(in_data_to_next_pe_16_25),
                        .Slide_data_26(in_data_to_next_pe_16_26), .Slide_data_27(in_data_to_next_pe_16_27),
                        .Slide_data_28(in_data_to_next_pe_16_28), .Slide_data_29(in_data_to_next_pe_16_29),
                        .Slide_data_30(in_data_to_next_pe_16_30), .Slide_data_31(in_data_to_next_pe_16_31),
                        .result(o_16),
                        .in_data_to_next_pe_0(in_data_to_next_pe_17_0), .in_data_to_next_pe_1(in_data_to_next_pe_17_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_17_2), .in_data_to_next_pe_3(in_data_to_next_pe_17_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_17_4), .in_data_to_next_pe_5(in_data_to_next_pe_17_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_17_6), .in_data_to_next_pe_7(in_data_to_next_pe_17_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_17_8), .in_data_to_next_pe_9(in_data_to_next_pe_17_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_17_10), .in_data_to_next_pe_11(in_data_to_next_pe_17_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_17_12), .in_data_to_next_pe_13(in_data_to_next_pe_17_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_17_14), .in_data_to_next_pe_15(in_data_to_next_pe_17_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_17_16), .in_data_to_next_pe_17(in_data_to_next_pe_17_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_17_18), .in_data_to_next_pe_19(in_data_to_next_pe_17_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_17_20), .in_data_to_next_pe_21(in_data_to_next_pe_17_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_17_22), .in_data_to_next_pe_23(in_data_to_next_pe_17_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_17_24), .in_data_to_next_pe_25(in_data_to_next_pe_17_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_17_26), .in_data_to_next_pe_27(in_data_to_next_pe_17_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_17_28), .in_data_to_next_pe_29(in_data_to_next_pe_17_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_17_30), .in_data_to_next_pe_31(in_data_to_next_pe_17_31),
                        .next_row_en(row_17_en)
        );
        
        PE_Row_B5   PE_R17_B5(   .clk(clk), .rst_n(row_17_en), .new_weight_val(new_weight_val[17]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_17_0), .Slide_data_1(in_data_to_next_pe_17_1),
                        .Slide_data_2(in_data_to_next_pe_17_2), .Slide_data_3(in_data_to_next_pe_17_3),
                        .Slide_data_4(in_data_to_next_pe_17_4), .Slide_data_5(in_data_to_next_pe_17_5),
                        .Slide_data_6(in_data_to_next_pe_17_6), .Slide_data_7(in_data_to_next_pe_17_7),
                        .Slide_data_8(in_data_to_next_pe_17_8), .Slide_data_9(in_data_to_next_pe_17_9),
                        .Slide_data_10(in_data_to_next_pe_17_10), .Slide_data_11(in_data_to_next_pe_17_11),
                        .Slide_data_12(in_data_to_next_pe_17_12), .Slide_data_13(in_data_to_next_pe_17_13),
                        .Slide_data_14(in_data_to_next_pe_17_14), .Slide_data_15(in_data_to_next_pe_17_15),
                        .Slide_data_16(in_data_to_next_pe_17_16), .Slide_data_17(in_data_to_next_pe_17_17),
                        .Slide_data_18(in_data_to_next_pe_17_18), .Slide_data_19(in_data_to_next_pe_17_19),
                        .Slide_data_20(in_data_to_next_pe_17_20), .Slide_data_21(in_data_to_next_pe_17_21),
                        .Slide_data_22(in_data_to_next_pe_17_22), .Slide_data_23(in_data_to_next_pe_17_23),
                        .Slide_data_24(in_data_to_next_pe_17_24), .Slide_data_25(in_data_to_next_pe_17_25),
                        .Slide_data_26(in_data_to_next_pe_17_26), .Slide_data_27(in_data_to_next_pe_17_27),
                        .Slide_data_28(in_data_to_next_pe_17_28), .Slide_data_29(in_data_to_next_pe_17_29),
                        .Slide_data_30(in_data_to_next_pe_17_30), .Slide_data_31(in_data_to_next_pe_17_31),
                        .result(o_17),
                        .in_data_to_next_pe_0(in_data_to_next_pe_18_0), .in_data_to_next_pe_1(in_data_to_next_pe_18_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_18_2), .in_data_to_next_pe_3(in_data_to_next_pe_18_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_18_4), .in_data_to_next_pe_5(in_data_to_next_pe_18_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_18_6), .in_data_to_next_pe_7(in_data_to_next_pe_18_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_18_8), .in_data_to_next_pe_9(in_data_to_next_pe_18_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_18_10), .in_data_to_next_pe_11(in_data_to_next_pe_18_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_18_12), .in_data_to_next_pe_13(in_data_to_next_pe_18_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_18_14), .in_data_to_next_pe_15(in_data_to_next_pe_18_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_18_16), .in_data_to_next_pe_17(in_data_to_next_pe_18_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_18_18), .in_data_to_next_pe_19(in_data_to_next_pe_18_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_18_20), .in_data_to_next_pe_21(in_data_to_next_pe_18_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_18_22), .in_data_to_next_pe_23(in_data_to_next_pe_18_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_18_24), .in_data_to_next_pe_25(in_data_to_next_pe_18_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_18_26), .in_data_to_next_pe_27(in_data_to_next_pe_18_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_18_28), .in_data_to_next_pe_29(in_data_to_next_pe_18_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_18_30), .in_data_to_next_pe_31(in_data_to_next_pe_18_31),
                        .next_row_en(row_18_en)
        );
        
        PE_Row_B5   PE_R18_B5(   .clk(clk), .rst_n(row_18_en), .new_weight_val(new_weight_val[18]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_18_0), .Slide_data_1(in_data_to_next_pe_18_1),
                        .Slide_data_2(in_data_to_next_pe_18_2), .Slide_data_3(in_data_to_next_pe_18_3),
                        .Slide_data_4(in_data_to_next_pe_18_4), .Slide_data_5(in_data_to_next_pe_18_5),
                        .Slide_data_6(in_data_to_next_pe_18_6), .Slide_data_7(in_data_to_next_pe_18_7),
                        .Slide_data_8(in_data_to_next_pe_18_8), .Slide_data_9(in_data_to_next_pe_18_9),
                        .Slide_data_10(in_data_to_next_pe_18_10), .Slide_data_11(in_data_to_next_pe_18_11),
                        .Slide_data_12(in_data_to_next_pe_18_12), .Slide_data_13(in_data_to_next_pe_18_13),
                        .Slide_data_14(in_data_to_next_pe_18_14), .Slide_data_15(in_data_to_next_pe_18_15),
                        .Slide_data_16(in_data_to_next_pe_18_16), .Slide_data_17(in_data_to_next_pe_18_17),
                        .Slide_data_18(in_data_to_next_pe_18_18), .Slide_data_19(in_data_to_next_pe_18_19),
                        .Slide_data_20(in_data_to_next_pe_18_20), .Slide_data_21(in_data_to_next_pe_18_21),
                        .Slide_data_22(in_data_to_next_pe_18_22), .Slide_data_23(in_data_to_next_pe_18_23),
                        .Slide_data_24(in_data_to_next_pe_18_24), .Slide_data_25(in_data_to_next_pe_18_25),
                        .Slide_data_26(in_data_to_next_pe_18_26), .Slide_data_27(in_data_to_next_pe_18_27),
                        .Slide_data_28(in_data_to_next_pe_18_28), .Slide_data_29(in_data_to_next_pe_18_29),
                        .Slide_data_30(in_data_to_next_pe_18_30), .Slide_data_31(in_data_to_next_pe_18_31),
                        .result(o_18),
                        .in_data_to_next_pe_0(in_data_to_next_pe_19_0), .in_data_to_next_pe_1(in_data_to_next_pe_19_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_19_2), .in_data_to_next_pe_3(in_data_to_next_pe_19_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_19_4), .in_data_to_next_pe_5(in_data_to_next_pe_19_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_19_6), .in_data_to_next_pe_7(in_data_to_next_pe_19_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_19_8), .in_data_to_next_pe_9(in_data_to_next_pe_19_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_19_10), .in_data_to_next_pe_11(in_data_to_next_pe_19_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_19_12), .in_data_to_next_pe_13(in_data_to_next_pe_19_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_19_14), .in_data_to_next_pe_15(in_data_to_next_pe_19_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_19_16), .in_data_to_next_pe_17(in_data_to_next_pe_19_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_19_18), .in_data_to_next_pe_19(in_data_to_next_pe_19_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_19_20), .in_data_to_next_pe_21(in_data_to_next_pe_19_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_19_22), .in_data_to_next_pe_23(in_data_to_next_pe_19_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_19_24), .in_data_to_next_pe_25(in_data_to_next_pe_19_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_19_26), .in_data_to_next_pe_27(in_data_to_next_pe_19_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_19_28), .in_data_to_next_pe_29(in_data_to_next_pe_19_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_19_30), .in_data_to_next_pe_31(in_data_to_next_pe_19_31),
                        .next_row_en(row_19_en)
        );
        
        PE_Row_B5   PE_R19_B5(   .clk(clk), .rst_n(row_19_en), .new_weight_val(new_weight_val[19]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_19_0), .Slide_data_1(in_data_to_next_pe_19_1),
                        .Slide_data_2(in_data_to_next_pe_19_2), .Slide_data_3(in_data_to_next_pe_19_3),
                        .Slide_data_4(in_data_to_next_pe_19_4), .Slide_data_5(in_data_to_next_pe_19_5),
                        .Slide_data_6(in_data_to_next_pe_19_6), .Slide_data_7(in_data_to_next_pe_19_7),
                        .Slide_data_8(in_data_to_next_pe_19_8), .Slide_data_9(in_data_to_next_pe_19_9),
                        .Slide_data_10(in_data_to_next_pe_19_10), .Slide_data_11(in_data_to_next_pe_19_11),
                        .Slide_data_12(in_data_to_next_pe_19_12), .Slide_data_13(in_data_to_next_pe_19_13),
                        .Slide_data_14(in_data_to_next_pe_19_14), .Slide_data_15(in_data_to_next_pe_19_15),
                        .Slide_data_16(in_data_to_next_pe_19_16), .Slide_data_17(in_data_to_next_pe_19_17),
                        .Slide_data_18(in_data_to_next_pe_19_18), .Slide_data_19(in_data_to_next_pe_19_19),
                        .Slide_data_20(in_data_to_next_pe_19_20), .Slide_data_21(in_data_to_next_pe_19_21),
                        .Slide_data_22(in_data_to_next_pe_19_22), .Slide_data_23(in_data_to_next_pe_19_23),
                        .Slide_data_24(in_data_to_next_pe_19_24), .Slide_data_25(in_data_to_next_pe_19_25),
                        .Slide_data_26(in_data_to_next_pe_19_26), .Slide_data_27(in_data_to_next_pe_19_27),
                        .Slide_data_28(in_data_to_next_pe_19_28), .Slide_data_29(in_data_to_next_pe_19_29),
                        .Slide_data_30(in_data_to_next_pe_19_30), .Slide_data_31(in_data_to_next_pe_19_31),
                        .result(o_19),
                        .in_data_to_next_pe_0(in_data_to_next_pe_20_0), .in_data_to_next_pe_1(in_data_to_next_pe_20_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_20_2), .in_data_to_next_pe_3(in_data_to_next_pe_20_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_20_4), .in_data_to_next_pe_5(in_data_to_next_pe_20_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_20_6), .in_data_to_next_pe_7(in_data_to_next_pe_20_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_20_8), .in_data_to_next_pe_9(in_data_to_next_pe_20_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_20_10), .in_data_to_next_pe_11(in_data_to_next_pe_20_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_20_12), .in_data_to_next_pe_13(in_data_to_next_pe_20_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_20_14), .in_data_to_next_pe_15(in_data_to_next_pe_20_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_20_16), .in_data_to_next_pe_17(in_data_to_next_pe_20_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_20_18), .in_data_to_next_pe_19(in_data_to_next_pe_20_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_20_20), .in_data_to_next_pe_21(in_data_to_next_pe_20_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_20_22), .in_data_to_next_pe_23(in_data_to_next_pe_20_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_20_24), .in_data_to_next_pe_25(in_data_to_next_pe_20_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_20_26), .in_data_to_next_pe_27(in_data_to_next_pe_20_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_20_28), .in_data_to_next_pe_29(in_data_to_next_pe_20_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_20_30), .in_data_to_next_pe_31(in_data_to_next_pe_20_31),
                        .next_row_en(row_20_en)
        );
        
        PE_Row_B5   PE_R20_B5(   .clk(clk), .rst_n(row_20_en), .new_weight_val(new_weight_val[20]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_20_0), .Slide_data_1(in_data_to_next_pe_20_1),
                        .Slide_data_2(in_data_to_next_pe_20_2), .Slide_data_3(in_data_to_next_pe_20_3),
                        .Slide_data_4(in_data_to_next_pe_20_4), .Slide_data_5(in_data_to_next_pe_20_5),
                        .Slide_data_6(in_data_to_next_pe_20_6), .Slide_data_7(in_data_to_next_pe_20_7),
                        .Slide_data_8(in_data_to_next_pe_20_8), .Slide_data_9(in_data_to_next_pe_20_9),
                        .Slide_data_10(in_data_to_next_pe_20_10), .Slide_data_11(in_data_to_next_pe_20_11),
                        .Slide_data_12(in_data_to_next_pe_20_12), .Slide_data_13(in_data_to_next_pe_20_13),
                        .Slide_data_14(in_data_to_next_pe_20_14), .Slide_data_15(in_data_to_next_pe_20_15),
                        .Slide_data_16(in_data_to_next_pe_20_16), .Slide_data_17(in_data_to_next_pe_20_17),
                        .Slide_data_18(in_data_to_next_pe_20_18), .Slide_data_19(in_data_to_next_pe_20_19),
                        .Slide_data_20(in_data_to_next_pe_20_20), .Slide_data_21(in_data_to_next_pe_20_21),
                        .Slide_data_22(in_data_to_next_pe_20_22), .Slide_data_23(in_data_to_next_pe_20_23),
                        .Slide_data_24(in_data_to_next_pe_20_24), .Slide_data_25(in_data_to_next_pe_20_25),
                        .Slide_data_26(in_data_to_next_pe_20_26), .Slide_data_27(in_data_to_next_pe_20_27),
                        .Slide_data_28(in_data_to_next_pe_20_28), .Slide_data_29(in_data_to_next_pe_20_29),
                        .Slide_data_30(in_data_to_next_pe_20_30), .Slide_data_31(in_data_to_next_pe_20_31),
                        .result(o_20),
                        .in_data_to_next_pe_0(in_data_to_next_pe_21_0), .in_data_to_next_pe_1(in_data_to_next_pe_21_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_21_2), .in_data_to_next_pe_3(in_data_to_next_pe_21_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_21_4), .in_data_to_next_pe_5(in_data_to_next_pe_21_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_21_6), .in_data_to_next_pe_7(in_data_to_next_pe_21_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_21_8), .in_data_to_next_pe_9(in_data_to_next_pe_21_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_21_10), .in_data_to_next_pe_11(in_data_to_next_pe_21_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_21_12), .in_data_to_next_pe_13(in_data_to_next_pe_21_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_21_14), .in_data_to_next_pe_15(in_data_to_next_pe_21_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_21_16), .in_data_to_next_pe_17(in_data_to_next_pe_21_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_21_18), .in_data_to_next_pe_19(in_data_to_next_pe_21_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_21_20), .in_data_to_next_pe_21(in_data_to_next_pe_21_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_21_22), .in_data_to_next_pe_23(in_data_to_next_pe_21_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_21_24), .in_data_to_next_pe_25(in_data_to_next_pe_21_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_21_26), .in_data_to_next_pe_27(in_data_to_next_pe_21_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_21_28), .in_data_to_next_pe_29(in_data_to_next_pe_21_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_21_30), .in_data_to_next_pe_31(in_data_to_next_pe_21_31),
                        .next_row_en(row_21_en)
        );
        
        PE_Row_B5   PE_R21_B5(   .clk(clk), .rst_n(row_21_en), .new_weight_val(new_weight_val[21]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_21_0), .Slide_data_1(in_data_to_next_pe_21_1),
                        .Slide_data_2(in_data_to_next_pe_21_2), .Slide_data_3(in_data_to_next_pe_21_3),
                        .Slide_data_4(in_data_to_next_pe_21_4), .Slide_data_5(in_data_to_next_pe_21_5),
                        .Slide_data_6(in_data_to_next_pe_21_6), .Slide_data_7(in_data_to_next_pe_21_7),
                        .Slide_data_8(in_data_to_next_pe_21_8), .Slide_data_9(in_data_to_next_pe_21_9),
                        .Slide_data_10(in_data_to_next_pe_21_10), .Slide_data_11(in_data_to_next_pe_21_11),
                        .Slide_data_12(in_data_to_next_pe_21_12), .Slide_data_13(in_data_to_next_pe_21_13),
                        .Slide_data_14(in_data_to_next_pe_21_14), .Slide_data_15(in_data_to_next_pe_21_15),
                        .Slide_data_16(in_data_to_next_pe_21_16), .Slide_data_17(in_data_to_next_pe_21_17),
                        .Slide_data_18(in_data_to_next_pe_21_18), .Slide_data_19(in_data_to_next_pe_21_19),
                        .Slide_data_20(in_data_to_next_pe_21_20), .Slide_data_21(in_data_to_next_pe_21_21),
                        .Slide_data_22(in_data_to_next_pe_21_22), .Slide_data_23(in_data_to_next_pe_21_23),
                        .Slide_data_24(in_data_to_next_pe_21_24), .Slide_data_25(in_data_to_next_pe_21_25),
                        .Slide_data_26(in_data_to_next_pe_21_26), .Slide_data_27(in_data_to_next_pe_21_27),
                        .Slide_data_28(in_data_to_next_pe_21_28), .Slide_data_29(in_data_to_next_pe_21_29),
                        .Slide_data_30(in_data_to_next_pe_21_30), .Slide_data_31(in_data_to_next_pe_21_31),
                        .result(o_21),
                        .in_data_to_next_pe_0(in_data_to_next_pe_22_0), .in_data_to_next_pe_1(in_data_to_next_pe_22_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_22_2), .in_data_to_next_pe_3(in_data_to_next_pe_22_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_22_4), .in_data_to_next_pe_5(in_data_to_next_pe_22_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_22_6), .in_data_to_next_pe_7(in_data_to_next_pe_22_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_22_8), .in_data_to_next_pe_9(in_data_to_next_pe_22_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_22_10), .in_data_to_next_pe_11(in_data_to_next_pe_22_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_22_12), .in_data_to_next_pe_13(in_data_to_next_pe_22_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_22_14), .in_data_to_next_pe_15(in_data_to_next_pe_22_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_22_16), .in_data_to_next_pe_17(in_data_to_next_pe_22_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_22_18), .in_data_to_next_pe_19(in_data_to_next_pe_22_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_22_20), .in_data_to_next_pe_21(in_data_to_next_pe_22_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_22_22), .in_data_to_next_pe_23(in_data_to_next_pe_22_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_22_24), .in_data_to_next_pe_25(in_data_to_next_pe_22_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_22_26), .in_data_to_next_pe_27(in_data_to_next_pe_22_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_22_28), .in_data_to_next_pe_29(in_data_to_next_pe_22_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_22_30), .in_data_to_next_pe_31(in_data_to_next_pe_22_31),
                        .next_row_en(row_22_en)
        );
        
        PE_Row_B5   PE_R22_B5(   .clk(clk), .rst_n(row_22_en), .new_weight_val(new_weight_val[22]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_22_0), .Slide_data_1(in_data_to_next_pe_22_1),
                        .Slide_data_2(in_data_to_next_pe_22_2), .Slide_data_3(in_data_to_next_pe_22_3),
                        .Slide_data_4(in_data_to_next_pe_22_4), .Slide_data_5(in_data_to_next_pe_22_5),
                        .Slide_data_6(in_data_to_next_pe_22_6), .Slide_data_7(in_data_to_next_pe_22_7),
                        .Slide_data_8(in_data_to_next_pe_22_8), .Slide_data_9(in_data_to_next_pe_22_9),
                        .Slide_data_10(in_data_to_next_pe_22_10), .Slide_data_11(in_data_to_next_pe_22_11),
                        .Slide_data_12(in_data_to_next_pe_22_12), .Slide_data_13(in_data_to_next_pe_22_13),
                        .Slide_data_14(in_data_to_next_pe_22_14), .Slide_data_15(in_data_to_next_pe_22_15),
                        .Slide_data_16(in_data_to_next_pe_22_16), .Slide_data_17(in_data_to_next_pe_22_17),
                        .Slide_data_18(in_data_to_next_pe_22_18), .Slide_data_19(in_data_to_next_pe_22_19),
                        .Slide_data_20(in_data_to_next_pe_22_20), .Slide_data_21(in_data_to_next_pe_22_21),
                        .Slide_data_22(in_data_to_next_pe_22_22), .Slide_data_23(in_data_to_next_pe_22_23),
                        .Slide_data_24(in_data_to_next_pe_22_24), .Slide_data_25(in_data_to_next_pe_22_25),
                        .Slide_data_26(in_data_to_next_pe_22_26), .Slide_data_27(in_data_to_next_pe_22_27),
                        .Slide_data_28(in_data_to_next_pe_22_28), .Slide_data_29(in_data_to_next_pe_22_29),
                        .Slide_data_30(in_data_to_next_pe_22_30), .Slide_data_31(in_data_to_next_pe_22_31),
                        .result(o_22),
                        .in_data_to_next_pe_0(in_data_to_next_pe_23_0), .in_data_to_next_pe_1(in_data_to_next_pe_23_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_23_2), .in_data_to_next_pe_3(in_data_to_next_pe_23_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_23_4), .in_data_to_next_pe_5(in_data_to_next_pe_23_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_23_6), .in_data_to_next_pe_7(in_data_to_next_pe_23_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_23_8), .in_data_to_next_pe_9(in_data_to_next_pe_23_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_23_10), .in_data_to_next_pe_11(in_data_to_next_pe_23_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_23_12), .in_data_to_next_pe_13(in_data_to_next_pe_23_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_23_14), .in_data_to_next_pe_15(in_data_to_next_pe_23_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_23_16), .in_data_to_next_pe_17(in_data_to_next_pe_23_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_23_18), .in_data_to_next_pe_19(in_data_to_next_pe_23_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_23_20), .in_data_to_next_pe_21(in_data_to_next_pe_23_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_23_22), .in_data_to_next_pe_23(in_data_to_next_pe_23_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_23_24), .in_data_to_next_pe_25(in_data_to_next_pe_23_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_23_26), .in_data_to_next_pe_27(in_data_to_next_pe_23_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_23_28), .in_data_to_next_pe_29(in_data_to_next_pe_23_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_23_30), .in_data_to_next_pe_31(in_data_to_next_pe_23_31),
                        .next_row_en(row_23_en)
        );
        
        PE_Row_B5   PE_R23_B5(   .clk(clk), .rst_n(row_23_en), .new_weight_val(new_weight_val[23]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_23_0), .Slide_data_1(in_data_to_next_pe_23_1),
                        .Slide_data_2(in_data_to_next_pe_23_2), .Slide_data_3(in_data_to_next_pe_23_3),
                        .Slide_data_4(in_data_to_next_pe_23_4), .Slide_data_5(in_data_to_next_pe_23_5),
                        .Slide_data_6(in_data_to_next_pe_23_6), .Slide_data_7(in_data_to_next_pe_23_7),
                        .Slide_data_8(in_data_to_next_pe_23_8), .Slide_data_9(in_data_to_next_pe_23_9),
                        .Slide_data_10(in_data_to_next_pe_23_10), .Slide_data_11(in_data_to_next_pe_23_11),
                        .Slide_data_12(in_data_to_next_pe_23_12), .Slide_data_13(in_data_to_next_pe_23_13),
                        .Slide_data_14(in_data_to_next_pe_23_14), .Slide_data_15(in_data_to_next_pe_23_15),
                        .Slide_data_16(in_data_to_next_pe_23_16), .Slide_data_17(in_data_to_next_pe_23_17),
                        .Slide_data_18(in_data_to_next_pe_23_18), .Slide_data_19(in_data_to_next_pe_23_19),
                        .Slide_data_20(in_data_to_next_pe_23_20), .Slide_data_21(in_data_to_next_pe_23_21),
                        .Slide_data_22(in_data_to_next_pe_23_22), .Slide_data_23(in_data_to_next_pe_23_23),
                        .Slide_data_24(in_data_to_next_pe_23_24), .Slide_data_25(in_data_to_next_pe_23_25),
                        .Slide_data_26(in_data_to_next_pe_23_26), .Slide_data_27(in_data_to_next_pe_23_27),
                        .Slide_data_28(in_data_to_next_pe_23_28), .Slide_data_29(in_data_to_next_pe_23_29),
                        .Slide_data_30(in_data_to_next_pe_23_30), .Slide_data_31(in_data_to_next_pe_23_31),
                        .result(o_23),
                        .in_data_to_next_pe_0(in_data_to_next_pe_24_0), .in_data_to_next_pe_1(in_data_to_next_pe_24_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_24_2), .in_data_to_next_pe_3(in_data_to_next_pe_24_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_24_4), .in_data_to_next_pe_5(in_data_to_next_pe_24_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_24_6), .in_data_to_next_pe_7(in_data_to_next_pe_24_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_24_8), .in_data_to_next_pe_9(in_data_to_next_pe_24_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_24_10), .in_data_to_next_pe_11(in_data_to_next_pe_24_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_24_12), .in_data_to_next_pe_13(in_data_to_next_pe_24_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_24_14), .in_data_to_next_pe_15(in_data_to_next_pe_24_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_24_16), .in_data_to_next_pe_17(in_data_to_next_pe_24_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_24_18), .in_data_to_next_pe_19(in_data_to_next_pe_24_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_24_20), .in_data_to_next_pe_21(in_data_to_next_pe_24_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_24_22), .in_data_to_next_pe_23(in_data_to_next_pe_24_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_24_24), .in_data_to_next_pe_25(in_data_to_next_pe_24_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_24_26), .in_data_to_next_pe_27(in_data_to_next_pe_24_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_24_28), .in_data_to_next_pe_29(in_data_to_next_pe_24_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_24_30), .in_data_to_next_pe_31(in_data_to_next_pe_24_31),
                        .next_row_en(row_24_en)
        );
        
        PE_Row_B5   PE_R24_B5(   .clk(clk), .rst_n(row_24_en), .new_weight_val(new_weight_val[24]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_24_0), .Slide_data_1(in_data_to_next_pe_24_1),
                        .Slide_data_2(in_data_to_next_pe_24_2), .Slide_data_3(in_data_to_next_pe_24_3),
                        .Slide_data_4(in_data_to_next_pe_24_4), .Slide_data_5(in_data_to_next_pe_24_5),
                        .Slide_data_6(in_data_to_next_pe_24_6), .Slide_data_7(in_data_to_next_pe_24_7),
                        .Slide_data_8(in_data_to_next_pe_24_8), .Slide_data_9(in_data_to_next_pe_24_9),
                        .Slide_data_10(in_data_to_next_pe_24_10), .Slide_data_11(in_data_to_next_pe_24_11),
                        .Slide_data_12(in_data_to_next_pe_24_12), .Slide_data_13(in_data_to_next_pe_24_13),
                        .Slide_data_14(in_data_to_next_pe_24_14), .Slide_data_15(in_data_to_next_pe_24_15),
                        .Slide_data_16(in_data_to_next_pe_24_16), .Slide_data_17(in_data_to_next_pe_24_17),
                        .Slide_data_18(in_data_to_next_pe_24_18), .Slide_data_19(in_data_to_next_pe_24_19),
                        .Slide_data_20(in_data_to_next_pe_24_20), .Slide_data_21(in_data_to_next_pe_24_21),
                        .Slide_data_22(in_data_to_next_pe_24_22), .Slide_data_23(in_data_to_next_pe_24_23),
                        .Slide_data_24(in_data_to_next_pe_24_24), .Slide_data_25(in_data_to_next_pe_24_25),
                        .Slide_data_26(in_data_to_next_pe_24_26), .Slide_data_27(in_data_to_next_pe_24_27),
                        .Slide_data_28(in_data_to_next_pe_24_28), .Slide_data_29(in_data_to_next_pe_24_29),
                        .Slide_data_30(in_data_to_next_pe_24_30), .Slide_data_31(in_data_to_next_pe_24_31),
                        .result(o_24),
                        .in_data_to_next_pe_0(in_data_to_next_pe_25_0), .in_data_to_next_pe_1(in_data_to_next_pe_25_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_25_2), .in_data_to_next_pe_3(in_data_to_next_pe_25_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_25_4), .in_data_to_next_pe_5(in_data_to_next_pe_25_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_25_6), .in_data_to_next_pe_7(in_data_to_next_pe_25_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_25_8), .in_data_to_next_pe_9(in_data_to_next_pe_25_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_25_10), .in_data_to_next_pe_11(in_data_to_next_pe_25_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_25_12), .in_data_to_next_pe_13(in_data_to_next_pe_25_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_25_14), .in_data_to_next_pe_15(in_data_to_next_pe_25_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_25_16), .in_data_to_next_pe_17(in_data_to_next_pe_25_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_25_18), .in_data_to_next_pe_19(in_data_to_next_pe_25_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_25_20), .in_data_to_next_pe_21(in_data_to_next_pe_25_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_25_22), .in_data_to_next_pe_23(in_data_to_next_pe_25_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_25_24), .in_data_to_next_pe_25(in_data_to_next_pe_25_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_25_26), .in_data_to_next_pe_27(in_data_to_next_pe_25_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_25_28), .in_data_to_next_pe_29(in_data_to_next_pe_25_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_25_30), .in_data_to_next_pe_31(in_data_to_next_pe_25_31),
                        .next_row_en(row_25_en)
        );
        
        PE_Row_B5   PE_R25_B5(   .clk(clk), .rst_n(row_25_en), .new_weight_val(new_weight_val[25]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_25_0), .Slide_data_1(in_data_to_next_pe_25_1),
                        .Slide_data_2(in_data_to_next_pe_25_2), .Slide_data_3(in_data_to_next_pe_25_3),
                        .Slide_data_4(in_data_to_next_pe_25_4), .Slide_data_5(in_data_to_next_pe_25_5),
                        .Slide_data_6(in_data_to_next_pe_25_6), .Slide_data_7(in_data_to_next_pe_25_7),
                        .Slide_data_8(in_data_to_next_pe_25_8), .Slide_data_9(in_data_to_next_pe_25_9),
                        .Slide_data_10(in_data_to_next_pe_25_10), .Slide_data_11(in_data_to_next_pe_25_11),
                        .Slide_data_12(in_data_to_next_pe_25_12), .Slide_data_13(in_data_to_next_pe_25_13),
                        .Slide_data_14(in_data_to_next_pe_25_14), .Slide_data_15(in_data_to_next_pe_25_15),
                        .Slide_data_16(in_data_to_next_pe_25_16), .Slide_data_17(in_data_to_next_pe_25_17),
                        .Slide_data_18(in_data_to_next_pe_25_18), .Slide_data_19(in_data_to_next_pe_25_19),
                        .Slide_data_20(in_data_to_next_pe_25_20), .Slide_data_21(in_data_to_next_pe_25_21),
                        .Slide_data_22(in_data_to_next_pe_25_22), .Slide_data_23(in_data_to_next_pe_25_23),
                        .Slide_data_24(in_data_to_next_pe_25_24), .Slide_data_25(in_data_to_next_pe_25_25),
                        .Slide_data_26(in_data_to_next_pe_25_26), .Slide_data_27(in_data_to_next_pe_25_27),
                        .Slide_data_28(in_data_to_next_pe_25_28), .Slide_data_29(in_data_to_next_pe_25_29),
                        .Slide_data_30(in_data_to_next_pe_25_30), .Slide_data_31(in_data_to_next_pe_25_31),
                        .result(o_25),
                        .in_data_to_next_pe_0(in_data_to_next_pe_26_0), .in_data_to_next_pe_1(in_data_to_next_pe_26_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_26_2), .in_data_to_next_pe_3(in_data_to_next_pe_26_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_26_4), .in_data_to_next_pe_5(in_data_to_next_pe_26_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_26_6), .in_data_to_next_pe_7(in_data_to_next_pe_26_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_26_8), .in_data_to_next_pe_9(in_data_to_next_pe_26_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_26_10), .in_data_to_next_pe_11(in_data_to_next_pe_26_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_26_12), .in_data_to_next_pe_13(in_data_to_next_pe_26_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_26_14), .in_data_to_next_pe_15(in_data_to_next_pe_26_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_26_16), .in_data_to_next_pe_17(in_data_to_next_pe_26_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_26_18), .in_data_to_next_pe_19(in_data_to_next_pe_26_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_26_20), .in_data_to_next_pe_21(in_data_to_next_pe_26_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_26_22), .in_data_to_next_pe_23(in_data_to_next_pe_26_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_26_24), .in_data_to_next_pe_25(in_data_to_next_pe_26_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_26_26), .in_data_to_next_pe_27(in_data_to_next_pe_26_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_26_28), .in_data_to_next_pe_29(in_data_to_next_pe_26_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_26_30), .in_data_to_next_pe_31(in_data_to_next_pe_26_31),
                        .next_row_en(row_26_en)
        );
        
        PE_Row_B5   PE_R26_B5(   .clk(clk), .rst_n(row_26_en), .new_weight_val(new_weight_val[26]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_26_0), .Slide_data_1(in_data_to_next_pe_26_1),
                        .Slide_data_2(in_data_to_next_pe_26_2), .Slide_data_3(in_data_to_next_pe_26_3),
                        .Slide_data_4(in_data_to_next_pe_26_4), .Slide_data_5(in_data_to_next_pe_26_5),
                        .Slide_data_6(in_data_to_next_pe_26_6), .Slide_data_7(in_data_to_next_pe_26_7),
                        .Slide_data_8(in_data_to_next_pe_26_8), .Slide_data_9(in_data_to_next_pe_26_9),
                        .Slide_data_10(in_data_to_next_pe_26_10), .Slide_data_11(in_data_to_next_pe_26_11),
                        .Slide_data_12(in_data_to_next_pe_26_12), .Slide_data_13(in_data_to_next_pe_26_13),
                        .Slide_data_14(in_data_to_next_pe_26_14), .Slide_data_15(in_data_to_next_pe_26_15),
                        .Slide_data_16(in_data_to_next_pe_26_16), .Slide_data_17(in_data_to_next_pe_26_17),
                        .Slide_data_18(in_data_to_next_pe_26_18), .Slide_data_19(in_data_to_next_pe_26_19),
                        .Slide_data_20(in_data_to_next_pe_26_20), .Slide_data_21(in_data_to_next_pe_26_21),
                        .Slide_data_22(in_data_to_next_pe_26_22), .Slide_data_23(in_data_to_next_pe_26_23),
                        .Slide_data_24(in_data_to_next_pe_26_24), .Slide_data_25(in_data_to_next_pe_26_25),
                        .Slide_data_26(in_data_to_next_pe_26_26), .Slide_data_27(in_data_to_next_pe_26_27),
                        .Slide_data_28(in_data_to_next_pe_26_28), .Slide_data_29(in_data_to_next_pe_26_29),
                        .Slide_data_30(in_data_to_next_pe_26_30), .Slide_data_31(in_data_to_next_pe_26_31),
                        .result(o_26),
                        .in_data_to_next_pe_0(in_data_to_next_pe_27_0), .in_data_to_next_pe_1(in_data_to_next_pe_27_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_27_2), .in_data_to_next_pe_3(in_data_to_next_pe_27_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_27_4), .in_data_to_next_pe_5(in_data_to_next_pe_27_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_27_6), .in_data_to_next_pe_7(in_data_to_next_pe_27_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_27_8), .in_data_to_next_pe_9(in_data_to_next_pe_27_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_27_10), .in_data_to_next_pe_11(in_data_to_next_pe_27_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_27_12), .in_data_to_next_pe_13(in_data_to_next_pe_27_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_27_14), .in_data_to_next_pe_15(in_data_to_next_pe_27_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_27_16), .in_data_to_next_pe_17(in_data_to_next_pe_27_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_27_18), .in_data_to_next_pe_19(in_data_to_next_pe_27_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_27_20), .in_data_to_next_pe_21(in_data_to_next_pe_27_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_27_22), .in_data_to_next_pe_23(in_data_to_next_pe_27_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_27_24), .in_data_to_next_pe_25(in_data_to_next_pe_27_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_27_26), .in_data_to_next_pe_27(in_data_to_next_pe_27_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_27_28), .in_data_to_next_pe_29(in_data_to_next_pe_27_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_27_30), .in_data_to_next_pe_31(in_data_to_next_pe_27_31),
                        .next_row_en(row_27_en)
        );
        
        PE_Row_B5   PE_R27_B5(   .clk(clk), .rst_n(row_27_en), .new_weight_val(new_weight_val[27]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_27_0), .Slide_data_1(in_data_to_next_pe_27_1),
                        .Slide_data_2(in_data_to_next_pe_27_2), .Slide_data_3(in_data_to_next_pe_27_3),
                        .Slide_data_4(in_data_to_next_pe_27_4), .Slide_data_5(in_data_to_next_pe_27_5),
                        .Slide_data_6(in_data_to_next_pe_27_6), .Slide_data_7(in_data_to_next_pe_27_7),
                        .Slide_data_8(in_data_to_next_pe_27_8), .Slide_data_9(in_data_to_next_pe_27_9),
                        .Slide_data_10(in_data_to_next_pe_27_10), .Slide_data_11(in_data_to_next_pe_27_11),
                        .Slide_data_12(in_data_to_next_pe_27_12), .Slide_data_13(in_data_to_next_pe_27_13),
                        .Slide_data_14(in_data_to_next_pe_27_14), .Slide_data_15(in_data_to_next_pe_27_15),
                        .Slide_data_16(in_data_to_next_pe_27_16), .Slide_data_17(in_data_to_next_pe_27_17),
                        .Slide_data_18(in_data_to_next_pe_27_18), .Slide_data_19(in_data_to_next_pe_27_19),
                        .Slide_data_20(in_data_to_next_pe_27_20), .Slide_data_21(in_data_to_next_pe_27_21),
                        .Slide_data_22(in_data_to_next_pe_27_22), .Slide_data_23(in_data_to_next_pe_27_23),
                        .Slide_data_24(in_data_to_next_pe_27_24), .Slide_data_25(in_data_to_next_pe_27_25),
                        .Slide_data_26(in_data_to_next_pe_27_26), .Slide_data_27(in_data_to_next_pe_27_27),
                        .Slide_data_28(in_data_to_next_pe_27_28), .Slide_data_29(in_data_to_next_pe_27_29),
                        .Slide_data_30(in_data_to_next_pe_27_30), .Slide_data_31(in_data_to_next_pe_27_31),
                        .result(o_27),
                        .in_data_to_next_pe_0(in_data_to_next_pe_28_0), .in_data_to_next_pe_1(in_data_to_next_pe_28_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_28_2), .in_data_to_next_pe_3(in_data_to_next_pe_28_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_28_4), .in_data_to_next_pe_5(in_data_to_next_pe_28_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_28_6), .in_data_to_next_pe_7(in_data_to_next_pe_28_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_28_8), .in_data_to_next_pe_9(in_data_to_next_pe_28_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_28_10), .in_data_to_next_pe_11(in_data_to_next_pe_28_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_28_12), .in_data_to_next_pe_13(in_data_to_next_pe_28_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_28_14), .in_data_to_next_pe_15(in_data_to_next_pe_28_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_28_16), .in_data_to_next_pe_17(in_data_to_next_pe_28_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_28_18), .in_data_to_next_pe_19(in_data_to_next_pe_28_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_28_20), .in_data_to_next_pe_21(in_data_to_next_pe_28_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_28_22), .in_data_to_next_pe_23(in_data_to_next_pe_28_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_28_24), .in_data_to_next_pe_25(in_data_to_next_pe_28_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_28_26), .in_data_to_next_pe_27(in_data_to_next_pe_28_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_28_28), .in_data_to_next_pe_29(in_data_to_next_pe_28_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_28_30), .in_data_to_next_pe_31(in_data_to_next_pe_28_31),
                        .next_row_en(row_28_en)
        );
        
        PE_Row_B5   PE_R28_B5(   .clk(clk), .rst_n(row_28_en), .new_weight_val(new_weight_val[28]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_28_0), .Slide_data_1(in_data_to_next_pe_28_1),
                        .Slide_data_2(in_data_to_next_pe_28_2), .Slide_data_3(in_data_to_next_pe_28_3),
                        .Slide_data_4(in_data_to_next_pe_28_4), .Slide_data_5(in_data_to_next_pe_28_5),
                        .Slide_data_6(in_data_to_next_pe_28_6), .Slide_data_7(in_data_to_next_pe_28_7),
                        .Slide_data_8(in_data_to_next_pe_28_8), .Slide_data_9(in_data_to_next_pe_28_9),
                        .Slide_data_10(in_data_to_next_pe_28_10), .Slide_data_11(in_data_to_next_pe_28_11),
                        .Slide_data_12(in_data_to_next_pe_28_12), .Slide_data_13(in_data_to_next_pe_28_13),
                        .Slide_data_14(in_data_to_next_pe_28_14), .Slide_data_15(in_data_to_next_pe_28_15),
                        .Slide_data_16(in_data_to_next_pe_28_16), .Slide_data_17(in_data_to_next_pe_28_17),
                        .Slide_data_18(in_data_to_next_pe_28_18), .Slide_data_19(in_data_to_next_pe_28_19),
                        .Slide_data_20(in_data_to_next_pe_28_20), .Slide_data_21(in_data_to_next_pe_28_21),
                        .Slide_data_22(in_data_to_next_pe_28_22), .Slide_data_23(in_data_to_next_pe_28_23),
                        .Slide_data_24(in_data_to_next_pe_28_24), .Slide_data_25(in_data_to_next_pe_28_25),
                        .Slide_data_26(in_data_to_next_pe_28_26), .Slide_data_27(in_data_to_next_pe_28_27),
                        .Slide_data_28(in_data_to_next_pe_28_28), .Slide_data_29(in_data_to_next_pe_28_29),
                        .Slide_data_30(in_data_to_next_pe_28_30), .Slide_data_31(in_data_to_next_pe_28_31),
                        .result(o_28),
                        .in_data_to_next_pe_0(in_data_to_next_pe_29_0), .in_data_to_next_pe_1(in_data_to_next_pe_29_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_29_2), .in_data_to_next_pe_3(in_data_to_next_pe_29_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_29_4), .in_data_to_next_pe_5(in_data_to_next_pe_29_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_29_6), .in_data_to_next_pe_7(in_data_to_next_pe_29_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_29_8), .in_data_to_next_pe_9(in_data_to_next_pe_29_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_29_10), .in_data_to_next_pe_11(in_data_to_next_pe_29_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_29_12), .in_data_to_next_pe_13(in_data_to_next_pe_29_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_29_14), .in_data_to_next_pe_15(in_data_to_next_pe_29_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_29_16), .in_data_to_next_pe_17(in_data_to_next_pe_29_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_29_18), .in_data_to_next_pe_19(in_data_to_next_pe_29_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_29_20), .in_data_to_next_pe_21(in_data_to_next_pe_29_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_29_22), .in_data_to_next_pe_23(in_data_to_next_pe_29_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_29_24), .in_data_to_next_pe_25(in_data_to_next_pe_29_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_29_26), .in_data_to_next_pe_27(in_data_to_next_pe_29_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_29_28), .in_data_to_next_pe_29(in_data_to_next_pe_29_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_29_30), .in_data_to_next_pe_31(in_data_to_next_pe_29_31),
                        .next_row_en(row_29_en)
        );
        
        PE_Row_B5   PE_R29_B5(   .clk(clk), .rst_n(row_29_en), .new_weight_val(new_weight_val[29]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_29_0), .Slide_data_1(in_data_to_next_pe_29_1),
                        .Slide_data_2(in_data_to_next_pe_29_2), .Slide_data_3(in_data_to_next_pe_29_3),
                        .Slide_data_4(in_data_to_next_pe_29_4), .Slide_data_5(in_data_to_next_pe_29_5),
                        .Slide_data_6(in_data_to_next_pe_29_6), .Slide_data_7(in_data_to_next_pe_29_7),
                        .Slide_data_8(in_data_to_next_pe_29_8), .Slide_data_9(in_data_to_next_pe_29_9),
                        .Slide_data_10(in_data_to_next_pe_29_10), .Slide_data_11(in_data_to_next_pe_29_11),
                        .Slide_data_12(in_data_to_next_pe_29_12), .Slide_data_13(in_data_to_next_pe_29_13),
                        .Slide_data_14(in_data_to_next_pe_29_14), .Slide_data_15(in_data_to_next_pe_29_15),
                        .Slide_data_16(in_data_to_next_pe_29_16), .Slide_data_17(in_data_to_next_pe_29_17),
                        .Slide_data_18(in_data_to_next_pe_29_18), .Slide_data_19(in_data_to_next_pe_29_19),
                        .Slide_data_20(in_data_to_next_pe_29_20), .Slide_data_21(in_data_to_next_pe_29_21),
                        .Slide_data_22(in_data_to_next_pe_29_22), .Slide_data_23(in_data_to_next_pe_29_23),
                        .Slide_data_24(in_data_to_next_pe_29_24), .Slide_data_25(in_data_to_next_pe_29_25),
                        .Slide_data_26(in_data_to_next_pe_29_26), .Slide_data_27(in_data_to_next_pe_29_27),
                        .Slide_data_28(in_data_to_next_pe_29_28), .Slide_data_29(in_data_to_next_pe_29_29),
                        .Slide_data_30(in_data_to_next_pe_29_30), .Slide_data_31(in_data_to_next_pe_29_31),
                        .result(o_29),
                        .in_data_to_next_pe_0(in_data_to_next_pe_30_0), .in_data_to_next_pe_1(in_data_to_next_pe_30_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_30_2), .in_data_to_next_pe_3(in_data_to_next_pe_30_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_30_4), .in_data_to_next_pe_5(in_data_to_next_pe_30_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_30_6), .in_data_to_next_pe_7(in_data_to_next_pe_30_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_30_8), .in_data_to_next_pe_9(in_data_to_next_pe_30_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_30_10), .in_data_to_next_pe_11(in_data_to_next_pe_30_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_30_12), .in_data_to_next_pe_13(in_data_to_next_pe_30_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_30_14), .in_data_to_next_pe_15(in_data_to_next_pe_30_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_30_16), .in_data_to_next_pe_17(in_data_to_next_pe_30_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_30_18), .in_data_to_next_pe_19(in_data_to_next_pe_30_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_30_20), .in_data_to_next_pe_21(in_data_to_next_pe_30_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_30_22), .in_data_to_next_pe_23(in_data_to_next_pe_30_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_30_24), .in_data_to_next_pe_25(in_data_to_next_pe_30_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_30_26), .in_data_to_next_pe_27(in_data_to_next_pe_30_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_30_28), .in_data_to_next_pe_29(in_data_to_next_pe_30_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_30_30), .in_data_to_next_pe_31(in_data_to_next_pe_30_31),
                        .next_row_en(row_30_en)
        );
        
        PE_Row_B5   PE_R30_B5(   .clk(clk), .rst_n(row_30_en), .new_weight_val(new_weight_val[30]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_30_0), .Slide_data_1(in_data_to_next_pe_30_1),
                        .Slide_data_2(in_data_to_next_pe_30_2), .Slide_data_3(in_data_to_next_pe_30_3),
                        .Slide_data_4(in_data_to_next_pe_30_4), .Slide_data_5(in_data_to_next_pe_30_5),
                        .Slide_data_6(in_data_to_next_pe_30_6), .Slide_data_7(in_data_to_next_pe_30_7),
                        .Slide_data_8(in_data_to_next_pe_30_8), .Slide_data_9(in_data_to_next_pe_30_9),
                        .Slide_data_10(in_data_to_next_pe_30_10), .Slide_data_11(in_data_to_next_pe_30_11),
                        .Slide_data_12(in_data_to_next_pe_30_12), .Slide_data_13(in_data_to_next_pe_30_13),
                        .Slide_data_14(in_data_to_next_pe_30_14), .Slide_data_15(in_data_to_next_pe_30_15),
                        .Slide_data_16(in_data_to_next_pe_30_16), .Slide_data_17(in_data_to_next_pe_30_17),
                        .Slide_data_18(in_data_to_next_pe_30_18), .Slide_data_19(in_data_to_next_pe_30_19),
                        .Slide_data_20(in_data_to_next_pe_30_20), .Slide_data_21(in_data_to_next_pe_30_21),
                        .Slide_data_22(in_data_to_next_pe_30_22), .Slide_data_23(in_data_to_next_pe_30_23),
                        .Slide_data_24(in_data_to_next_pe_30_24), .Slide_data_25(in_data_to_next_pe_30_25),
                        .Slide_data_26(in_data_to_next_pe_30_26), .Slide_data_27(in_data_to_next_pe_30_27),
                        .Slide_data_28(in_data_to_next_pe_30_28), .Slide_data_29(in_data_to_next_pe_30_29),
                        .Slide_data_30(in_data_to_next_pe_30_30), .Slide_data_31(in_data_to_next_pe_30_31),
                        .result(o_30),
                        .in_data_to_next_pe_0(in_data_to_next_pe_31_0), .in_data_to_next_pe_1(in_data_to_next_pe_31_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_31_2), .in_data_to_next_pe_3(in_data_to_next_pe_31_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_31_4), .in_data_to_next_pe_5(in_data_to_next_pe_31_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_31_6), .in_data_to_next_pe_7(in_data_to_next_pe_31_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_31_8), .in_data_to_next_pe_9(in_data_to_next_pe_31_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_31_10), .in_data_to_next_pe_11(in_data_to_next_pe_31_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_31_12), .in_data_to_next_pe_13(in_data_to_next_pe_31_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_31_14), .in_data_to_next_pe_15(in_data_to_next_pe_31_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_31_16), .in_data_to_next_pe_17(in_data_to_next_pe_31_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_31_18), .in_data_to_next_pe_19(in_data_to_next_pe_31_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_31_20), .in_data_to_next_pe_21(in_data_to_next_pe_31_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_31_22), .in_data_to_next_pe_23(in_data_to_next_pe_31_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_31_24), .in_data_to_next_pe_25(in_data_to_next_pe_31_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_31_26), .in_data_to_next_pe_27(in_data_to_next_pe_31_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_31_28), .in_data_to_next_pe_29(in_data_to_next_pe_31_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_31_30), .in_data_to_next_pe_31(in_data_to_next_pe_31_31),
                        .next_row_en(row_31_en)
        );
        
        PE_Row_B5   PE_R31_B5(   .clk(clk), .rst_n(row_31_en), .new_weight_val(new_weight_val[31]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_31_0), .Slide_data_1(in_data_to_next_pe_31_1),
                        .Slide_data_2(in_data_to_next_pe_31_2), .Slide_data_3(in_data_to_next_pe_31_3),
                        .Slide_data_4(in_data_to_next_pe_31_4), .Slide_data_5(in_data_to_next_pe_31_5),
                        .Slide_data_6(in_data_to_next_pe_31_6), .Slide_data_7(in_data_to_next_pe_31_7),
                        .Slide_data_8(in_data_to_next_pe_31_8), .Slide_data_9(in_data_to_next_pe_31_9),
                        .Slide_data_10(in_data_to_next_pe_31_10), .Slide_data_11(in_data_to_next_pe_31_11),
                        .Slide_data_12(in_data_to_next_pe_31_12), .Slide_data_13(in_data_to_next_pe_31_13),
                        .Slide_data_14(in_data_to_next_pe_31_14), .Slide_data_15(in_data_to_next_pe_31_15),
                        .Slide_data_16(in_data_to_next_pe_31_16), .Slide_data_17(in_data_to_next_pe_31_17),
                        .Slide_data_18(in_data_to_next_pe_31_18), .Slide_data_19(in_data_to_next_pe_31_19),
                        .Slide_data_20(in_data_to_next_pe_31_20), .Slide_data_21(in_data_to_next_pe_31_21),
                        .Slide_data_22(in_data_to_next_pe_31_22), .Slide_data_23(in_data_to_next_pe_31_23),
                        .Slide_data_24(in_data_to_next_pe_31_24), .Slide_data_25(in_data_to_next_pe_31_25),
                        .Slide_data_26(in_data_to_next_pe_31_26), .Slide_data_27(in_data_to_next_pe_31_27),
                        .Slide_data_28(in_data_to_next_pe_31_28), .Slide_data_29(in_data_to_next_pe_31_29),
                        .Slide_data_30(in_data_to_next_pe_31_30), .Slide_data_31(in_data_to_next_pe_31_31),
                        .result(o_31),
                        .in_data_to_next_pe_0(in_data_to_next_pe_32_0), .in_data_to_next_pe_1(in_data_to_next_pe_32_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_32_2), .in_data_to_next_pe_3(in_data_to_next_pe_32_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_32_4), .in_data_to_next_pe_5(in_data_to_next_pe_32_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_32_6), .in_data_to_next_pe_7(in_data_to_next_pe_32_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_32_8), .in_data_to_next_pe_9(in_data_to_next_pe_32_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_32_10), .in_data_to_next_pe_11(in_data_to_next_pe_32_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_32_12), .in_data_to_next_pe_13(in_data_to_next_pe_32_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_32_14), .in_data_to_next_pe_15(in_data_to_next_pe_32_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_32_16), .in_data_to_next_pe_17(in_data_to_next_pe_32_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_32_18), .in_data_to_next_pe_19(in_data_to_next_pe_32_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_32_20), .in_data_to_next_pe_21(in_data_to_next_pe_32_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_32_22), .in_data_to_next_pe_23(in_data_to_next_pe_32_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_32_24), .in_data_to_next_pe_25(in_data_to_next_pe_32_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_32_26), .in_data_to_next_pe_27(in_data_to_next_pe_32_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_32_28), .in_data_to_next_pe_29(in_data_to_next_pe_32_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_32_30), .in_data_to_next_pe_31(in_data_to_next_pe_32_31),
                        .next_row_en(row_32_en)
        );
        
        PE_Row_B5   PE_R32_B5(   .clk(clk), .rst_n(row_32_en), .new_weight_val(new_weight_val[32]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_32_0), .Slide_data_1(in_data_to_next_pe_32_1),
                        .Slide_data_2(in_data_to_next_pe_32_2), .Slide_data_3(in_data_to_next_pe_32_3),
                        .Slide_data_4(in_data_to_next_pe_32_4), .Slide_data_5(in_data_to_next_pe_32_5),
                        .Slide_data_6(in_data_to_next_pe_32_6), .Slide_data_7(in_data_to_next_pe_32_7),
                        .Slide_data_8(in_data_to_next_pe_32_8), .Slide_data_9(in_data_to_next_pe_32_9),
                        .Slide_data_10(in_data_to_next_pe_32_10), .Slide_data_11(in_data_to_next_pe_32_11),
                        .Slide_data_12(in_data_to_next_pe_32_12), .Slide_data_13(in_data_to_next_pe_32_13),
                        .Slide_data_14(in_data_to_next_pe_32_14), .Slide_data_15(in_data_to_next_pe_32_15),
                        .Slide_data_16(in_data_to_next_pe_32_16), .Slide_data_17(in_data_to_next_pe_32_17),
                        .Slide_data_18(in_data_to_next_pe_32_18), .Slide_data_19(in_data_to_next_pe_32_19),
                        .Slide_data_20(in_data_to_next_pe_32_20), .Slide_data_21(in_data_to_next_pe_32_21),
                        .Slide_data_22(in_data_to_next_pe_32_22), .Slide_data_23(in_data_to_next_pe_32_23),
                        .Slide_data_24(in_data_to_next_pe_32_24), .Slide_data_25(in_data_to_next_pe_32_25),
                        .Slide_data_26(in_data_to_next_pe_32_26), .Slide_data_27(in_data_to_next_pe_32_27),
                        .Slide_data_28(in_data_to_next_pe_32_28), .Slide_data_29(in_data_to_next_pe_32_29),
                        .Slide_data_30(in_data_to_next_pe_32_30), .Slide_data_31(in_data_to_next_pe_32_31),
                        .result(o_32),
                        .in_data_to_next_pe_0(in_data_to_next_pe_33_0), .in_data_to_next_pe_1(in_data_to_next_pe_33_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_33_2), .in_data_to_next_pe_3(in_data_to_next_pe_33_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_33_4), .in_data_to_next_pe_5(in_data_to_next_pe_33_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_33_6), .in_data_to_next_pe_7(in_data_to_next_pe_33_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_33_8), .in_data_to_next_pe_9(in_data_to_next_pe_33_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_33_10), .in_data_to_next_pe_11(in_data_to_next_pe_33_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_33_12), .in_data_to_next_pe_13(in_data_to_next_pe_33_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_33_14), .in_data_to_next_pe_15(in_data_to_next_pe_33_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_33_16), .in_data_to_next_pe_17(in_data_to_next_pe_33_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_33_18), .in_data_to_next_pe_19(in_data_to_next_pe_33_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_33_20), .in_data_to_next_pe_21(in_data_to_next_pe_33_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_33_22), .in_data_to_next_pe_23(in_data_to_next_pe_33_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_33_24), .in_data_to_next_pe_25(in_data_to_next_pe_33_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_33_26), .in_data_to_next_pe_27(in_data_to_next_pe_33_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_33_28), .in_data_to_next_pe_29(in_data_to_next_pe_33_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_33_30), .in_data_to_next_pe_31(in_data_to_next_pe_33_31),
                        .next_row_en(row_33_en)
        );
        
        PE_Row_B5   PE_R33_B5(   .clk(clk), .rst_n(row_33_en), .new_weight_val(new_weight_val[33]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_33_0), .Slide_data_1(in_data_to_next_pe_33_1),
                        .Slide_data_2(in_data_to_next_pe_33_2), .Slide_data_3(in_data_to_next_pe_33_3),
                        .Slide_data_4(in_data_to_next_pe_33_4), .Slide_data_5(in_data_to_next_pe_33_5),
                        .Slide_data_6(in_data_to_next_pe_33_6), .Slide_data_7(in_data_to_next_pe_33_7),
                        .Slide_data_8(in_data_to_next_pe_33_8), .Slide_data_9(in_data_to_next_pe_33_9),
                        .Slide_data_10(in_data_to_next_pe_33_10), .Slide_data_11(in_data_to_next_pe_33_11),
                        .Slide_data_12(in_data_to_next_pe_33_12), .Slide_data_13(in_data_to_next_pe_33_13),
                        .Slide_data_14(in_data_to_next_pe_33_14), .Slide_data_15(in_data_to_next_pe_33_15),
                        .Slide_data_16(in_data_to_next_pe_33_16), .Slide_data_17(in_data_to_next_pe_33_17),
                        .Slide_data_18(in_data_to_next_pe_33_18), .Slide_data_19(in_data_to_next_pe_33_19),
                        .Slide_data_20(in_data_to_next_pe_33_20), .Slide_data_21(in_data_to_next_pe_33_21),
                        .Slide_data_22(in_data_to_next_pe_33_22), .Slide_data_23(in_data_to_next_pe_33_23),
                        .Slide_data_24(in_data_to_next_pe_33_24), .Slide_data_25(in_data_to_next_pe_33_25),
                        .Slide_data_26(in_data_to_next_pe_33_26), .Slide_data_27(in_data_to_next_pe_33_27),
                        .Slide_data_28(in_data_to_next_pe_33_28), .Slide_data_29(in_data_to_next_pe_33_29),
                        .Slide_data_30(in_data_to_next_pe_33_30), .Slide_data_31(in_data_to_next_pe_33_31),
                        .result(o_33),
                        .in_data_to_next_pe_0(in_data_to_next_pe_34_0), .in_data_to_next_pe_1(in_data_to_next_pe_34_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_34_2), .in_data_to_next_pe_3(in_data_to_next_pe_34_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_34_4), .in_data_to_next_pe_5(in_data_to_next_pe_34_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_34_6), .in_data_to_next_pe_7(in_data_to_next_pe_34_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_34_8), .in_data_to_next_pe_9(in_data_to_next_pe_34_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_34_10), .in_data_to_next_pe_11(in_data_to_next_pe_34_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_34_12), .in_data_to_next_pe_13(in_data_to_next_pe_34_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_34_14), .in_data_to_next_pe_15(in_data_to_next_pe_34_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_34_16), .in_data_to_next_pe_17(in_data_to_next_pe_34_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_34_18), .in_data_to_next_pe_19(in_data_to_next_pe_34_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_34_20), .in_data_to_next_pe_21(in_data_to_next_pe_34_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_34_22), .in_data_to_next_pe_23(in_data_to_next_pe_34_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_34_24), .in_data_to_next_pe_25(in_data_to_next_pe_34_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_34_26), .in_data_to_next_pe_27(in_data_to_next_pe_34_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_34_28), .in_data_to_next_pe_29(in_data_to_next_pe_34_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_34_30), .in_data_to_next_pe_31(in_data_to_next_pe_34_31),
                        .next_row_en(row_34_en)
        );
        
        PE_Row_B5   PE_R34_B5(   .clk(clk), .rst_n(row_34_en), .new_weight_val(new_weight_val[34]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_34_0), .Slide_data_1(in_data_to_next_pe_34_1),
                        .Slide_data_2(in_data_to_next_pe_34_2), .Slide_data_3(in_data_to_next_pe_34_3),
                        .Slide_data_4(in_data_to_next_pe_34_4), .Slide_data_5(in_data_to_next_pe_34_5),
                        .Slide_data_6(in_data_to_next_pe_34_6), .Slide_data_7(in_data_to_next_pe_34_7),
                        .Slide_data_8(in_data_to_next_pe_34_8), .Slide_data_9(in_data_to_next_pe_34_9),
                        .Slide_data_10(in_data_to_next_pe_34_10), .Slide_data_11(in_data_to_next_pe_34_11),
                        .Slide_data_12(in_data_to_next_pe_34_12), .Slide_data_13(in_data_to_next_pe_34_13),
                        .Slide_data_14(in_data_to_next_pe_34_14), .Slide_data_15(in_data_to_next_pe_34_15),
                        .Slide_data_16(in_data_to_next_pe_34_16), .Slide_data_17(in_data_to_next_pe_34_17),
                        .Slide_data_18(in_data_to_next_pe_34_18), .Slide_data_19(in_data_to_next_pe_34_19),
                        .Slide_data_20(in_data_to_next_pe_34_20), .Slide_data_21(in_data_to_next_pe_34_21),
                        .Slide_data_22(in_data_to_next_pe_34_22), .Slide_data_23(in_data_to_next_pe_34_23),
                        .Slide_data_24(in_data_to_next_pe_34_24), .Slide_data_25(in_data_to_next_pe_34_25),
                        .Slide_data_26(in_data_to_next_pe_34_26), .Slide_data_27(in_data_to_next_pe_34_27),
                        .Slide_data_28(in_data_to_next_pe_34_28), .Slide_data_29(in_data_to_next_pe_34_29),
                        .Slide_data_30(in_data_to_next_pe_34_30), .Slide_data_31(in_data_to_next_pe_34_31),
                        .result(o_34),
                        .in_data_to_next_pe_0(in_data_to_next_pe_35_0), .in_data_to_next_pe_1(in_data_to_next_pe_35_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_35_2), .in_data_to_next_pe_3(in_data_to_next_pe_35_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_35_4), .in_data_to_next_pe_5(in_data_to_next_pe_35_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_35_6), .in_data_to_next_pe_7(in_data_to_next_pe_35_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_35_8), .in_data_to_next_pe_9(in_data_to_next_pe_35_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_35_10), .in_data_to_next_pe_11(in_data_to_next_pe_35_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_35_12), .in_data_to_next_pe_13(in_data_to_next_pe_35_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_35_14), .in_data_to_next_pe_15(in_data_to_next_pe_35_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_35_16), .in_data_to_next_pe_17(in_data_to_next_pe_35_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_35_18), .in_data_to_next_pe_19(in_data_to_next_pe_35_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_35_20), .in_data_to_next_pe_21(in_data_to_next_pe_35_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_35_22), .in_data_to_next_pe_23(in_data_to_next_pe_35_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_35_24), .in_data_to_next_pe_25(in_data_to_next_pe_35_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_35_26), .in_data_to_next_pe_27(in_data_to_next_pe_35_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_35_28), .in_data_to_next_pe_29(in_data_to_next_pe_35_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_35_30), .in_data_to_next_pe_31(in_data_to_next_pe_35_31),
                        .next_row_en(row_35_en)
        );
        
        PE_Row_B5   PE_R35_B5(   .clk(clk), .rst_n(row_35_en), .new_weight_val(new_weight_val[35]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_35_0), .Slide_data_1(in_data_to_next_pe_35_1),
                        .Slide_data_2(in_data_to_next_pe_35_2), .Slide_data_3(in_data_to_next_pe_35_3),
                        .Slide_data_4(in_data_to_next_pe_35_4), .Slide_data_5(in_data_to_next_pe_35_5),
                        .Slide_data_6(in_data_to_next_pe_35_6), .Slide_data_7(in_data_to_next_pe_35_7),
                        .Slide_data_8(in_data_to_next_pe_35_8), .Slide_data_9(in_data_to_next_pe_35_9),
                        .Slide_data_10(in_data_to_next_pe_35_10), .Slide_data_11(in_data_to_next_pe_35_11),
                        .Slide_data_12(in_data_to_next_pe_35_12), .Slide_data_13(in_data_to_next_pe_35_13),
                        .Slide_data_14(in_data_to_next_pe_35_14), .Slide_data_15(in_data_to_next_pe_35_15),
                        .Slide_data_16(in_data_to_next_pe_35_16), .Slide_data_17(in_data_to_next_pe_35_17),
                        .Slide_data_18(in_data_to_next_pe_35_18), .Slide_data_19(in_data_to_next_pe_35_19),
                        .Slide_data_20(in_data_to_next_pe_35_20), .Slide_data_21(in_data_to_next_pe_35_21),
                        .Slide_data_22(in_data_to_next_pe_35_22), .Slide_data_23(in_data_to_next_pe_35_23),
                        .Slide_data_24(in_data_to_next_pe_35_24), .Slide_data_25(in_data_to_next_pe_35_25),
                        .Slide_data_26(in_data_to_next_pe_35_26), .Slide_data_27(in_data_to_next_pe_35_27),
                        .Slide_data_28(in_data_to_next_pe_35_28), .Slide_data_29(in_data_to_next_pe_35_29),
                        .Slide_data_30(in_data_to_next_pe_35_30), .Slide_data_31(in_data_to_next_pe_35_31),
                        .result(o_35),
                        .in_data_to_next_pe_0(in_data_to_next_pe_36_0), .in_data_to_next_pe_1(in_data_to_next_pe_36_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_36_2), .in_data_to_next_pe_3(in_data_to_next_pe_36_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_36_4), .in_data_to_next_pe_5(in_data_to_next_pe_36_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_36_6), .in_data_to_next_pe_7(in_data_to_next_pe_36_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_36_8), .in_data_to_next_pe_9(in_data_to_next_pe_36_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_36_10), .in_data_to_next_pe_11(in_data_to_next_pe_36_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_36_12), .in_data_to_next_pe_13(in_data_to_next_pe_36_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_36_14), .in_data_to_next_pe_15(in_data_to_next_pe_36_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_36_16), .in_data_to_next_pe_17(in_data_to_next_pe_36_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_36_18), .in_data_to_next_pe_19(in_data_to_next_pe_36_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_36_20), .in_data_to_next_pe_21(in_data_to_next_pe_36_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_36_22), .in_data_to_next_pe_23(in_data_to_next_pe_36_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_36_24), .in_data_to_next_pe_25(in_data_to_next_pe_36_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_36_26), .in_data_to_next_pe_27(in_data_to_next_pe_36_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_36_28), .in_data_to_next_pe_29(in_data_to_next_pe_36_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_36_30), .in_data_to_next_pe_31(in_data_to_next_pe_36_31),
                        .next_row_en(row_36_en)
        );
        
        PE_Row_B5   PE_R36_B5(   .clk(clk), .rst_n(row_36_en), .new_weight_val(new_weight_val[36]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_36_0), .Slide_data_1(in_data_to_next_pe_36_1),
                        .Slide_data_2(in_data_to_next_pe_36_2), .Slide_data_3(in_data_to_next_pe_36_3),
                        .Slide_data_4(in_data_to_next_pe_36_4), .Slide_data_5(in_data_to_next_pe_36_5),
                        .Slide_data_6(in_data_to_next_pe_36_6), .Slide_data_7(in_data_to_next_pe_36_7),
                        .Slide_data_8(in_data_to_next_pe_36_8), .Slide_data_9(in_data_to_next_pe_36_9),
                        .Slide_data_10(in_data_to_next_pe_36_10), .Slide_data_11(in_data_to_next_pe_36_11),
                        .Slide_data_12(in_data_to_next_pe_36_12), .Slide_data_13(in_data_to_next_pe_36_13),
                        .Slide_data_14(in_data_to_next_pe_36_14), .Slide_data_15(in_data_to_next_pe_36_15),
                        .Slide_data_16(in_data_to_next_pe_36_16), .Slide_data_17(in_data_to_next_pe_36_17),
                        .Slide_data_18(in_data_to_next_pe_36_18), .Slide_data_19(in_data_to_next_pe_36_19),
                        .Slide_data_20(in_data_to_next_pe_36_20), .Slide_data_21(in_data_to_next_pe_36_21),
                        .Slide_data_22(in_data_to_next_pe_36_22), .Slide_data_23(in_data_to_next_pe_36_23),
                        .Slide_data_24(in_data_to_next_pe_36_24), .Slide_data_25(in_data_to_next_pe_36_25),
                        .Slide_data_26(in_data_to_next_pe_36_26), .Slide_data_27(in_data_to_next_pe_36_27),
                        .Slide_data_28(in_data_to_next_pe_36_28), .Slide_data_29(in_data_to_next_pe_36_29),
                        .Slide_data_30(in_data_to_next_pe_36_30), .Slide_data_31(in_data_to_next_pe_36_31),
                        .result(o_36),
                        .in_data_to_next_pe_0(in_data_to_next_pe_37_0), .in_data_to_next_pe_1(in_data_to_next_pe_37_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_37_2), .in_data_to_next_pe_3(in_data_to_next_pe_37_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_37_4), .in_data_to_next_pe_5(in_data_to_next_pe_37_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_37_6), .in_data_to_next_pe_7(in_data_to_next_pe_37_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_37_8), .in_data_to_next_pe_9(in_data_to_next_pe_37_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_37_10), .in_data_to_next_pe_11(in_data_to_next_pe_37_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_37_12), .in_data_to_next_pe_13(in_data_to_next_pe_37_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_37_14), .in_data_to_next_pe_15(in_data_to_next_pe_37_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_37_16), .in_data_to_next_pe_17(in_data_to_next_pe_37_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_37_18), .in_data_to_next_pe_19(in_data_to_next_pe_37_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_37_20), .in_data_to_next_pe_21(in_data_to_next_pe_37_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_37_22), .in_data_to_next_pe_23(in_data_to_next_pe_37_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_37_24), .in_data_to_next_pe_25(in_data_to_next_pe_37_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_37_26), .in_data_to_next_pe_27(in_data_to_next_pe_37_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_37_28), .in_data_to_next_pe_29(in_data_to_next_pe_37_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_37_30), .in_data_to_next_pe_31(in_data_to_next_pe_37_31),
                        .next_row_en(row_37_en)
        );
        
        PE_Row_B5   PE_R37_B5(   .clk(clk), .rst_n(row_37_en), .new_weight_val(new_weight_val[37]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_37_0), .Slide_data_1(in_data_to_next_pe_37_1),
                        .Slide_data_2(in_data_to_next_pe_37_2), .Slide_data_3(in_data_to_next_pe_37_3),
                        .Slide_data_4(in_data_to_next_pe_37_4), .Slide_data_5(in_data_to_next_pe_37_5),
                        .Slide_data_6(in_data_to_next_pe_37_6), .Slide_data_7(in_data_to_next_pe_37_7),
                        .Slide_data_8(in_data_to_next_pe_37_8), .Slide_data_9(in_data_to_next_pe_37_9),
                        .Slide_data_10(in_data_to_next_pe_37_10), .Slide_data_11(in_data_to_next_pe_37_11),
                        .Slide_data_12(in_data_to_next_pe_37_12), .Slide_data_13(in_data_to_next_pe_37_13),
                        .Slide_data_14(in_data_to_next_pe_37_14), .Slide_data_15(in_data_to_next_pe_37_15),
                        .Slide_data_16(in_data_to_next_pe_37_16), .Slide_data_17(in_data_to_next_pe_37_17),
                        .Slide_data_18(in_data_to_next_pe_37_18), .Slide_data_19(in_data_to_next_pe_37_19),
                        .Slide_data_20(in_data_to_next_pe_37_20), .Slide_data_21(in_data_to_next_pe_37_21),
                        .Slide_data_22(in_data_to_next_pe_37_22), .Slide_data_23(in_data_to_next_pe_37_23),
                        .Slide_data_24(in_data_to_next_pe_37_24), .Slide_data_25(in_data_to_next_pe_37_25),
                        .Slide_data_26(in_data_to_next_pe_37_26), .Slide_data_27(in_data_to_next_pe_37_27),
                        .Slide_data_28(in_data_to_next_pe_37_28), .Slide_data_29(in_data_to_next_pe_37_29),
                        .Slide_data_30(in_data_to_next_pe_37_30), .Slide_data_31(in_data_to_next_pe_37_31),
                        .result(o_37),
                        .in_data_to_next_pe_0(in_data_to_next_pe_38_0), .in_data_to_next_pe_1(in_data_to_next_pe_38_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_38_2), .in_data_to_next_pe_3(in_data_to_next_pe_38_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_38_4), .in_data_to_next_pe_5(in_data_to_next_pe_38_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_38_6), .in_data_to_next_pe_7(in_data_to_next_pe_38_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_38_8), .in_data_to_next_pe_9(in_data_to_next_pe_38_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_38_10), .in_data_to_next_pe_11(in_data_to_next_pe_38_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_38_12), .in_data_to_next_pe_13(in_data_to_next_pe_38_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_38_14), .in_data_to_next_pe_15(in_data_to_next_pe_38_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_38_16), .in_data_to_next_pe_17(in_data_to_next_pe_38_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_38_18), .in_data_to_next_pe_19(in_data_to_next_pe_38_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_38_20), .in_data_to_next_pe_21(in_data_to_next_pe_38_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_38_22), .in_data_to_next_pe_23(in_data_to_next_pe_38_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_38_24), .in_data_to_next_pe_25(in_data_to_next_pe_38_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_38_26), .in_data_to_next_pe_27(in_data_to_next_pe_38_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_38_28), .in_data_to_next_pe_29(in_data_to_next_pe_38_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_38_30), .in_data_to_next_pe_31(in_data_to_next_pe_38_31),
                        .next_row_en(row_38_en)
        );
        
        PE_Row_B5   PE_R38_B5(   .clk(clk), .rst_n(row_38_en), .new_weight_val(new_weight_val[38]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_38_0), .Slide_data_1(in_data_to_next_pe_38_1),
                        .Slide_data_2(in_data_to_next_pe_38_2), .Slide_data_3(in_data_to_next_pe_38_3),
                        .Slide_data_4(in_data_to_next_pe_38_4), .Slide_data_5(in_data_to_next_pe_38_5),
                        .Slide_data_6(in_data_to_next_pe_38_6), .Slide_data_7(in_data_to_next_pe_38_7),
                        .Slide_data_8(in_data_to_next_pe_38_8), .Slide_data_9(in_data_to_next_pe_38_9),
                        .Slide_data_10(in_data_to_next_pe_38_10), .Slide_data_11(in_data_to_next_pe_38_11),
                        .Slide_data_12(in_data_to_next_pe_38_12), .Slide_data_13(in_data_to_next_pe_38_13),
                        .Slide_data_14(in_data_to_next_pe_38_14), .Slide_data_15(in_data_to_next_pe_38_15),
                        .Slide_data_16(in_data_to_next_pe_38_16), .Slide_data_17(in_data_to_next_pe_38_17),
                        .Slide_data_18(in_data_to_next_pe_38_18), .Slide_data_19(in_data_to_next_pe_38_19),
                        .Slide_data_20(in_data_to_next_pe_38_20), .Slide_data_21(in_data_to_next_pe_38_21),
                        .Slide_data_22(in_data_to_next_pe_38_22), .Slide_data_23(in_data_to_next_pe_38_23),
                        .Slide_data_24(in_data_to_next_pe_38_24), .Slide_data_25(in_data_to_next_pe_38_25),
                        .Slide_data_26(in_data_to_next_pe_38_26), .Slide_data_27(in_data_to_next_pe_38_27),
                        .Slide_data_28(in_data_to_next_pe_38_28), .Slide_data_29(in_data_to_next_pe_38_29),
                        .Slide_data_30(in_data_to_next_pe_38_30), .Slide_data_31(in_data_to_next_pe_38_31),
                        .result(o_38),
                        .in_data_to_next_pe_0(in_data_to_next_pe_39_0), .in_data_to_next_pe_1(in_data_to_next_pe_39_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_39_2), .in_data_to_next_pe_3(in_data_to_next_pe_39_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_39_4), .in_data_to_next_pe_5(in_data_to_next_pe_39_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_39_6), .in_data_to_next_pe_7(in_data_to_next_pe_39_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_39_8), .in_data_to_next_pe_9(in_data_to_next_pe_39_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_39_10), .in_data_to_next_pe_11(in_data_to_next_pe_39_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_39_12), .in_data_to_next_pe_13(in_data_to_next_pe_39_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_39_14), .in_data_to_next_pe_15(in_data_to_next_pe_39_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_39_16), .in_data_to_next_pe_17(in_data_to_next_pe_39_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_39_18), .in_data_to_next_pe_19(in_data_to_next_pe_39_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_39_20), .in_data_to_next_pe_21(in_data_to_next_pe_39_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_39_22), .in_data_to_next_pe_23(in_data_to_next_pe_39_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_39_24), .in_data_to_next_pe_25(in_data_to_next_pe_39_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_39_26), .in_data_to_next_pe_27(in_data_to_next_pe_39_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_39_28), .in_data_to_next_pe_29(in_data_to_next_pe_39_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_39_30), .in_data_to_next_pe_31(in_data_to_next_pe_39_31),
                        .next_row_en(row_39_en)
        );
        
        PE_Row_B5   PE_R39_B5(   .clk(clk), .rst_n(row_39_en), .new_weight_val(new_weight_val[39]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_39_0), .Slide_data_1(in_data_to_next_pe_39_1),
                        .Slide_data_2(in_data_to_next_pe_39_2), .Slide_data_3(in_data_to_next_pe_39_3),
                        .Slide_data_4(in_data_to_next_pe_39_4), .Slide_data_5(in_data_to_next_pe_39_5),
                        .Slide_data_6(in_data_to_next_pe_39_6), .Slide_data_7(in_data_to_next_pe_39_7),
                        .Slide_data_8(in_data_to_next_pe_39_8), .Slide_data_9(in_data_to_next_pe_39_9),
                        .Slide_data_10(in_data_to_next_pe_39_10), .Slide_data_11(in_data_to_next_pe_39_11),
                        .Slide_data_12(in_data_to_next_pe_39_12), .Slide_data_13(in_data_to_next_pe_39_13),
                        .Slide_data_14(in_data_to_next_pe_39_14), .Slide_data_15(in_data_to_next_pe_39_15),
                        .Slide_data_16(in_data_to_next_pe_39_16), .Slide_data_17(in_data_to_next_pe_39_17),
                        .Slide_data_18(in_data_to_next_pe_39_18), .Slide_data_19(in_data_to_next_pe_39_19),
                        .Slide_data_20(in_data_to_next_pe_39_20), .Slide_data_21(in_data_to_next_pe_39_21),
                        .Slide_data_22(in_data_to_next_pe_39_22), .Slide_data_23(in_data_to_next_pe_39_23),
                        .Slide_data_24(in_data_to_next_pe_39_24), .Slide_data_25(in_data_to_next_pe_39_25),
                        .Slide_data_26(in_data_to_next_pe_39_26), .Slide_data_27(in_data_to_next_pe_39_27),
                        .Slide_data_28(in_data_to_next_pe_39_28), .Slide_data_29(in_data_to_next_pe_39_29),
                        .Slide_data_30(in_data_to_next_pe_39_30), .Slide_data_31(in_data_to_next_pe_39_31),
                        .result(o_39),
                        .in_data_to_next_pe_0(in_data_to_next_pe_40_0), .in_data_to_next_pe_1(in_data_to_next_pe_40_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_40_2), .in_data_to_next_pe_3(in_data_to_next_pe_40_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_40_4), .in_data_to_next_pe_5(in_data_to_next_pe_40_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_40_6), .in_data_to_next_pe_7(in_data_to_next_pe_40_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_40_8), .in_data_to_next_pe_9(in_data_to_next_pe_40_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_40_10), .in_data_to_next_pe_11(in_data_to_next_pe_40_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_40_12), .in_data_to_next_pe_13(in_data_to_next_pe_40_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_40_14), .in_data_to_next_pe_15(in_data_to_next_pe_40_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_40_16), .in_data_to_next_pe_17(in_data_to_next_pe_40_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_40_18), .in_data_to_next_pe_19(in_data_to_next_pe_40_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_40_20), .in_data_to_next_pe_21(in_data_to_next_pe_40_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_40_22), .in_data_to_next_pe_23(in_data_to_next_pe_40_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_40_24), .in_data_to_next_pe_25(in_data_to_next_pe_40_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_40_26), .in_data_to_next_pe_27(in_data_to_next_pe_40_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_40_28), .in_data_to_next_pe_29(in_data_to_next_pe_40_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_40_30), .in_data_to_next_pe_31(in_data_to_next_pe_40_31),
                        .next_row_en(row_40_en)
        );
        
        PE_Row_B5   PE_R40_B5(   .clk(clk), .rst_n(row_40_en), .new_weight_val(new_weight_val[40]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_40_0), .Slide_data_1(in_data_to_next_pe_40_1),
                        .Slide_data_2(in_data_to_next_pe_40_2), .Slide_data_3(in_data_to_next_pe_40_3),
                        .Slide_data_4(in_data_to_next_pe_40_4), .Slide_data_5(in_data_to_next_pe_40_5),
                        .Slide_data_6(in_data_to_next_pe_40_6), .Slide_data_7(in_data_to_next_pe_40_7),
                        .Slide_data_8(in_data_to_next_pe_40_8), .Slide_data_9(in_data_to_next_pe_40_9),
                        .Slide_data_10(in_data_to_next_pe_40_10), .Slide_data_11(in_data_to_next_pe_40_11),
                        .Slide_data_12(in_data_to_next_pe_40_12), .Slide_data_13(in_data_to_next_pe_40_13),
                        .Slide_data_14(in_data_to_next_pe_40_14), .Slide_data_15(in_data_to_next_pe_40_15),
                        .Slide_data_16(in_data_to_next_pe_40_16), .Slide_data_17(in_data_to_next_pe_40_17),
                        .Slide_data_18(in_data_to_next_pe_40_18), .Slide_data_19(in_data_to_next_pe_40_19),
                        .Slide_data_20(in_data_to_next_pe_40_20), .Slide_data_21(in_data_to_next_pe_40_21),
                        .Slide_data_22(in_data_to_next_pe_40_22), .Slide_data_23(in_data_to_next_pe_40_23),
                        .Slide_data_24(in_data_to_next_pe_40_24), .Slide_data_25(in_data_to_next_pe_40_25),
                        .Slide_data_26(in_data_to_next_pe_40_26), .Slide_data_27(in_data_to_next_pe_40_27),
                        .Slide_data_28(in_data_to_next_pe_40_28), .Slide_data_29(in_data_to_next_pe_40_29),
                        .Slide_data_30(in_data_to_next_pe_40_30), .Slide_data_31(in_data_to_next_pe_40_31),
                        .result(o_40),
                        .in_data_to_next_pe_0(in_data_to_next_pe_41_0), .in_data_to_next_pe_1(in_data_to_next_pe_41_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_41_2), .in_data_to_next_pe_3(in_data_to_next_pe_41_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_41_4), .in_data_to_next_pe_5(in_data_to_next_pe_41_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_41_6), .in_data_to_next_pe_7(in_data_to_next_pe_41_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_41_8), .in_data_to_next_pe_9(in_data_to_next_pe_41_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_41_10), .in_data_to_next_pe_11(in_data_to_next_pe_41_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_41_12), .in_data_to_next_pe_13(in_data_to_next_pe_41_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_41_14), .in_data_to_next_pe_15(in_data_to_next_pe_41_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_41_16), .in_data_to_next_pe_17(in_data_to_next_pe_41_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_41_18), .in_data_to_next_pe_19(in_data_to_next_pe_41_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_41_20), .in_data_to_next_pe_21(in_data_to_next_pe_41_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_41_22), .in_data_to_next_pe_23(in_data_to_next_pe_41_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_41_24), .in_data_to_next_pe_25(in_data_to_next_pe_41_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_41_26), .in_data_to_next_pe_27(in_data_to_next_pe_41_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_41_28), .in_data_to_next_pe_29(in_data_to_next_pe_41_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_41_30), .in_data_to_next_pe_31(in_data_to_next_pe_41_31),
                        .next_row_en(row_41_en)
        );
        
        PE_Row_B5   PE_R41_B5(   .clk(clk), .rst_n(row_41_en), .new_weight_val(new_weight_val[41]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_41_0), .Slide_data_1(in_data_to_next_pe_41_1),
                        .Slide_data_2(in_data_to_next_pe_41_2), .Slide_data_3(in_data_to_next_pe_41_3),
                        .Slide_data_4(in_data_to_next_pe_41_4), .Slide_data_5(in_data_to_next_pe_41_5),
                        .Slide_data_6(in_data_to_next_pe_41_6), .Slide_data_7(in_data_to_next_pe_41_7),
                        .Slide_data_8(in_data_to_next_pe_41_8), .Slide_data_9(in_data_to_next_pe_41_9),
                        .Slide_data_10(in_data_to_next_pe_41_10), .Slide_data_11(in_data_to_next_pe_41_11),
                        .Slide_data_12(in_data_to_next_pe_41_12), .Slide_data_13(in_data_to_next_pe_41_13),
                        .Slide_data_14(in_data_to_next_pe_41_14), .Slide_data_15(in_data_to_next_pe_41_15),
                        .Slide_data_16(in_data_to_next_pe_41_16), .Slide_data_17(in_data_to_next_pe_41_17),
                        .Slide_data_18(in_data_to_next_pe_41_18), .Slide_data_19(in_data_to_next_pe_41_19),
                        .Slide_data_20(in_data_to_next_pe_41_20), .Slide_data_21(in_data_to_next_pe_41_21),
                        .Slide_data_22(in_data_to_next_pe_41_22), .Slide_data_23(in_data_to_next_pe_41_23),
                        .Slide_data_24(in_data_to_next_pe_41_24), .Slide_data_25(in_data_to_next_pe_41_25),
                        .Slide_data_26(in_data_to_next_pe_41_26), .Slide_data_27(in_data_to_next_pe_41_27),
                        .Slide_data_28(in_data_to_next_pe_41_28), .Slide_data_29(in_data_to_next_pe_41_29),
                        .Slide_data_30(in_data_to_next_pe_41_30), .Slide_data_31(in_data_to_next_pe_41_31),
                        .result(o_41),
                        .in_data_to_next_pe_0(in_data_to_next_pe_42_0), .in_data_to_next_pe_1(in_data_to_next_pe_42_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_42_2), .in_data_to_next_pe_3(in_data_to_next_pe_42_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_42_4), .in_data_to_next_pe_5(in_data_to_next_pe_42_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_42_6), .in_data_to_next_pe_7(in_data_to_next_pe_42_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_42_8), .in_data_to_next_pe_9(in_data_to_next_pe_42_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_42_10), .in_data_to_next_pe_11(in_data_to_next_pe_42_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_42_12), .in_data_to_next_pe_13(in_data_to_next_pe_42_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_42_14), .in_data_to_next_pe_15(in_data_to_next_pe_42_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_42_16), .in_data_to_next_pe_17(in_data_to_next_pe_42_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_42_18), .in_data_to_next_pe_19(in_data_to_next_pe_42_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_42_20), .in_data_to_next_pe_21(in_data_to_next_pe_42_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_42_22), .in_data_to_next_pe_23(in_data_to_next_pe_42_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_42_24), .in_data_to_next_pe_25(in_data_to_next_pe_42_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_42_26), .in_data_to_next_pe_27(in_data_to_next_pe_42_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_42_28), .in_data_to_next_pe_29(in_data_to_next_pe_42_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_42_30), .in_data_to_next_pe_31(in_data_to_next_pe_42_31),
                        .next_row_en(row_42_en)
        );
        
        PE_Row_B5   PE_R42_B5(   .clk(clk), .rst_n(row_42_en), .new_weight_val(new_weight_val[42]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_42_0), .Slide_data_1(in_data_to_next_pe_42_1),
                        .Slide_data_2(in_data_to_next_pe_42_2), .Slide_data_3(in_data_to_next_pe_42_3),
                        .Slide_data_4(in_data_to_next_pe_42_4), .Slide_data_5(in_data_to_next_pe_42_5),
                        .Slide_data_6(in_data_to_next_pe_42_6), .Slide_data_7(in_data_to_next_pe_42_7),
                        .Slide_data_8(in_data_to_next_pe_42_8), .Slide_data_9(in_data_to_next_pe_42_9),
                        .Slide_data_10(in_data_to_next_pe_42_10), .Slide_data_11(in_data_to_next_pe_42_11),
                        .Slide_data_12(in_data_to_next_pe_42_12), .Slide_data_13(in_data_to_next_pe_42_13),
                        .Slide_data_14(in_data_to_next_pe_42_14), .Slide_data_15(in_data_to_next_pe_42_15),
                        .Slide_data_16(in_data_to_next_pe_42_16), .Slide_data_17(in_data_to_next_pe_42_17),
                        .Slide_data_18(in_data_to_next_pe_42_18), .Slide_data_19(in_data_to_next_pe_42_19),
                        .Slide_data_20(in_data_to_next_pe_42_20), .Slide_data_21(in_data_to_next_pe_42_21),
                        .Slide_data_22(in_data_to_next_pe_42_22), .Slide_data_23(in_data_to_next_pe_42_23),
                        .Slide_data_24(in_data_to_next_pe_42_24), .Slide_data_25(in_data_to_next_pe_42_25),
                        .Slide_data_26(in_data_to_next_pe_42_26), .Slide_data_27(in_data_to_next_pe_42_27),
                        .Slide_data_28(in_data_to_next_pe_42_28), .Slide_data_29(in_data_to_next_pe_42_29),
                        .Slide_data_30(in_data_to_next_pe_42_30), .Slide_data_31(in_data_to_next_pe_42_31),
                        .result(o_42),
                        .in_data_to_next_pe_0(in_data_to_next_pe_43_0), .in_data_to_next_pe_1(in_data_to_next_pe_43_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_43_2), .in_data_to_next_pe_3(in_data_to_next_pe_43_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_43_4), .in_data_to_next_pe_5(in_data_to_next_pe_43_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_43_6), .in_data_to_next_pe_7(in_data_to_next_pe_43_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_43_8), .in_data_to_next_pe_9(in_data_to_next_pe_43_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_43_10), .in_data_to_next_pe_11(in_data_to_next_pe_43_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_43_12), .in_data_to_next_pe_13(in_data_to_next_pe_43_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_43_14), .in_data_to_next_pe_15(in_data_to_next_pe_43_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_43_16), .in_data_to_next_pe_17(in_data_to_next_pe_43_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_43_18), .in_data_to_next_pe_19(in_data_to_next_pe_43_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_43_20), .in_data_to_next_pe_21(in_data_to_next_pe_43_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_43_22), .in_data_to_next_pe_23(in_data_to_next_pe_43_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_43_24), .in_data_to_next_pe_25(in_data_to_next_pe_43_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_43_26), .in_data_to_next_pe_27(in_data_to_next_pe_43_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_43_28), .in_data_to_next_pe_29(in_data_to_next_pe_43_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_43_30), .in_data_to_next_pe_31(in_data_to_next_pe_43_31),
                        .next_row_en(row_43_en)
        );
        
        PE_Row_B5   PE_R43_B5(   .clk(clk), .rst_n(row_43_en), .new_weight_val(new_weight_val[43]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_43_0), .Slide_data_1(in_data_to_next_pe_43_1),
                        .Slide_data_2(in_data_to_next_pe_43_2), .Slide_data_3(in_data_to_next_pe_43_3),
                        .Slide_data_4(in_data_to_next_pe_43_4), .Slide_data_5(in_data_to_next_pe_43_5),
                        .Slide_data_6(in_data_to_next_pe_43_6), .Slide_data_7(in_data_to_next_pe_43_7),
                        .Slide_data_8(in_data_to_next_pe_43_8), .Slide_data_9(in_data_to_next_pe_43_9),
                        .Slide_data_10(in_data_to_next_pe_43_10), .Slide_data_11(in_data_to_next_pe_43_11),
                        .Slide_data_12(in_data_to_next_pe_43_12), .Slide_data_13(in_data_to_next_pe_43_13),
                        .Slide_data_14(in_data_to_next_pe_43_14), .Slide_data_15(in_data_to_next_pe_43_15),
                        .Slide_data_16(in_data_to_next_pe_43_16), .Slide_data_17(in_data_to_next_pe_43_17),
                        .Slide_data_18(in_data_to_next_pe_43_18), .Slide_data_19(in_data_to_next_pe_43_19),
                        .Slide_data_20(in_data_to_next_pe_43_20), .Slide_data_21(in_data_to_next_pe_43_21),
                        .Slide_data_22(in_data_to_next_pe_43_22), .Slide_data_23(in_data_to_next_pe_43_23),
                        .Slide_data_24(in_data_to_next_pe_43_24), .Slide_data_25(in_data_to_next_pe_43_25),
                        .Slide_data_26(in_data_to_next_pe_43_26), .Slide_data_27(in_data_to_next_pe_43_27),
                        .Slide_data_28(in_data_to_next_pe_43_28), .Slide_data_29(in_data_to_next_pe_43_29),
                        .Slide_data_30(in_data_to_next_pe_43_30), .Slide_data_31(in_data_to_next_pe_43_31),
                        .result(o_43),
                        .in_data_to_next_pe_0(in_data_to_next_pe_44_0), .in_data_to_next_pe_1(in_data_to_next_pe_44_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_44_2), .in_data_to_next_pe_3(in_data_to_next_pe_44_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_44_4), .in_data_to_next_pe_5(in_data_to_next_pe_44_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_44_6), .in_data_to_next_pe_7(in_data_to_next_pe_44_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_44_8), .in_data_to_next_pe_9(in_data_to_next_pe_44_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_44_10), .in_data_to_next_pe_11(in_data_to_next_pe_44_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_44_12), .in_data_to_next_pe_13(in_data_to_next_pe_44_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_44_14), .in_data_to_next_pe_15(in_data_to_next_pe_44_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_44_16), .in_data_to_next_pe_17(in_data_to_next_pe_44_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_44_18), .in_data_to_next_pe_19(in_data_to_next_pe_44_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_44_20), .in_data_to_next_pe_21(in_data_to_next_pe_44_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_44_22), .in_data_to_next_pe_23(in_data_to_next_pe_44_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_44_24), .in_data_to_next_pe_25(in_data_to_next_pe_44_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_44_26), .in_data_to_next_pe_27(in_data_to_next_pe_44_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_44_28), .in_data_to_next_pe_29(in_data_to_next_pe_44_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_44_30), .in_data_to_next_pe_31(in_data_to_next_pe_44_31),
                        .next_row_en(row_44_en)
        );
        
        PE_Row_B5   PE_R44_B5(   .clk(clk), .rst_n(row_44_en), .new_weight_val(new_weight_val[44]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_44_0), .Slide_data_1(in_data_to_next_pe_44_1),
                        .Slide_data_2(in_data_to_next_pe_44_2), .Slide_data_3(in_data_to_next_pe_44_3),
                        .Slide_data_4(in_data_to_next_pe_44_4), .Slide_data_5(in_data_to_next_pe_44_5),
                        .Slide_data_6(in_data_to_next_pe_44_6), .Slide_data_7(in_data_to_next_pe_44_7),
                        .Slide_data_8(in_data_to_next_pe_44_8), .Slide_data_9(in_data_to_next_pe_44_9),
                        .Slide_data_10(in_data_to_next_pe_44_10), .Slide_data_11(in_data_to_next_pe_44_11),
                        .Slide_data_12(in_data_to_next_pe_44_12), .Slide_data_13(in_data_to_next_pe_44_13),
                        .Slide_data_14(in_data_to_next_pe_44_14), .Slide_data_15(in_data_to_next_pe_44_15),
                        .Slide_data_16(in_data_to_next_pe_44_16), .Slide_data_17(in_data_to_next_pe_44_17),
                        .Slide_data_18(in_data_to_next_pe_44_18), .Slide_data_19(in_data_to_next_pe_44_19),
                        .Slide_data_20(in_data_to_next_pe_44_20), .Slide_data_21(in_data_to_next_pe_44_21),
                        .Slide_data_22(in_data_to_next_pe_44_22), .Slide_data_23(in_data_to_next_pe_44_23),
                        .Slide_data_24(in_data_to_next_pe_44_24), .Slide_data_25(in_data_to_next_pe_44_25),
                        .Slide_data_26(in_data_to_next_pe_44_26), .Slide_data_27(in_data_to_next_pe_44_27),
                        .Slide_data_28(in_data_to_next_pe_44_28), .Slide_data_29(in_data_to_next_pe_44_29),
                        .Slide_data_30(in_data_to_next_pe_44_30), .Slide_data_31(in_data_to_next_pe_44_31),
                        .result(o_44),
                        .in_data_to_next_pe_0(in_data_to_next_pe_45_0), .in_data_to_next_pe_1(in_data_to_next_pe_45_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_45_2), .in_data_to_next_pe_3(in_data_to_next_pe_45_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_45_4), .in_data_to_next_pe_5(in_data_to_next_pe_45_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_45_6), .in_data_to_next_pe_7(in_data_to_next_pe_45_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_45_8), .in_data_to_next_pe_9(in_data_to_next_pe_45_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_45_10), .in_data_to_next_pe_11(in_data_to_next_pe_45_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_45_12), .in_data_to_next_pe_13(in_data_to_next_pe_45_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_45_14), .in_data_to_next_pe_15(in_data_to_next_pe_45_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_45_16), .in_data_to_next_pe_17(in_data_to_next_pe_45_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_45_18), .in_data_to_next_pe_19(in_data_to_next_pe_45_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_45_20), .in_data_to_next_pe_21(in_data_to_next_pe_45_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_45_22), .in_data_to_next_pe_23(in_data_to_next_pe_45_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_45_24), .in_data_to_next_pe_25(in_data_to_next_pe_45_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_45_26), .in_data_to_next_pe_27(in_data_to_next_pe_45_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_45_28), .in_data_to_next_pe_29(in_data_to_next_pe_45_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_45_30), .in_data_to_next_pe_31(in_data_to_next_pe_45_31),
                        .next_row_en(row_45_en)
        );
        
        PE_Row_B5   PE_R45_B5(   .clk(clk), .rst_n(row_45_en), .new_weight_val(new_weight_val[45]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_45_0), .Slide_data_1(in_data_to_next_pe_45_1),
                        .Slide_data_2(in_data_to_next_pe_45_2), .Slide_data_3(in_data_to_next_pe_45_3),
                        .Slide_data_4(in_data_to_next_pe_45_4), .Slide_data_5(in_data_to_next_pe_45_5),
                        .Slide_data_6(in_data_to_next_pe_45_6), .Slide_data_7(in_data_to_next_pe_45_7),
                        .Slide_data_8(in_data_to_next_pe_45_8), .Slide_data_9(in_data_to_next_pe_45_9),
                        .Slide_data_10(in_data_to_next_pe_45_10), .Slide_data_11(in_data_to_next_pe_45_11),
                        .Slide_data_12(in_data_to_next_pe_45_12), .Slide_data_13(in_data_to_next_pe_45_13),
                        .Slide_data_14(in_data_to_next_pe_45_14), .Slide_data_15(in_data_to_next_pe_45_15),
                        .Slide_data_16(in_data_to_next_pe_45_16), .Slide_data_17(in_data_to_next_pe_45_17),
                        .Slide_data_18(in_data_to_next_pe_45_18), .Slide_data_19(in_data_to_next_pe_45_19),
                        .Slide_data_20(in_data_to_next_pe_45_20), .Slide_data_21(in_data_to_next_pe_45_21),
                        .Slide_data_22(in_data_to_next_pe_45_22), .Slide_data_23(in_data_to_next_pe_45_23),
                        .Slide_data_24(in_data_to_next_pe_45_24), .Slide_data_25(in_data_to_next_pe_45_25),
                        .Slide_data_26(in_data_to_next_pe_45_26), .Slide_data_27(in_data_to_next_pe_45_27),
                        .Slide_data_28(in_data_to_next_pe_45_28), .Slide_data_29(in_data_to_next_pe_45_29),
                        .Slide_data_30(in_data_to_next_pe_45_30), .Slide_data_31(in_data_to_next_pe_45_31),
                        .result(o_45),
                        .in_data_to_next_pe_0(in_data_to_next_pe_46_0), .in_data_to_next_pe_1(in_data_to_next_pe_46_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_46_2), .in_data_to_next_pe_3(in_data_to_next_pe_46_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_46_4), .in_data_to_next_pe_5(in_data_to_next_pe_46_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_46_6), .in_data_to_next_pe_7(in_data_to_next_pe_46_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_46_8), .in_data_to_next_pe_9(in_data_to_next_pe_46_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_46_10), .in_data_to_next_pe_11(in_data_to_next_pe_46_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_46_12), .in_data_to_next_pe_13(in_data_to_next_pe_46_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_46_14), .in_data_to_next_pe_15(in_data_to_next_pe_46_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_46_16), .in_data_to_next_pe_17(in_data_to_next_pe_46_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_46_18), .in_data_to_next_pe_19(in_data_to_next_pe_46_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_46_20), .in_data_to_next_pe_21(in_data_to_next_pe_46_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_46_22), .in_data_to_next_pe_23(in_data_to_next_pe_46_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_46_24), .in_data_to_next_pe_25(in_data_to_next_pe_46_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_46_26), .in_data_to_next_pe_27(in_data_to_next_pe_46_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_46_28), .in_data_to_next_pe_29(in_data_to_next_pe_46_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_46_30), .in_data_to_next_pe_31(in_data_to_next_pe_46_31),
                        .next_row_en(row_46_en)
        );
        
        PE_Row_B5   PE_R46_B5(   .clk(clk), .rst_n(row_46_en), .new_weight_val(new_weight_val[46]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_46_0), .Slide_data_1(in_data_to_next_pe_46_1),
                        .Slide_data_2(in_data_to_next_pe_46_2), .Slide_data_3(in_data_to_next_pe_46_3),
                        .Slide_data_4(in_data_to_next_pe_46_4), .Slide_data_5(in_data_to_next_pe_46_5),
                        .Slide_data_6(in_data_to_next_pe_46_6), .Slide_data_7(in_data_to_next_pe_46_7),
                        .Slide_data_8(in_data_to_next_pe_46_8), .Slide_data_9(in_data_to_next_pe_46_9),
                        .Slide_data_10(in_data_to_next_pe_46_10), .Slide_data_11(in_data_to_next_pe_46_11),
                        .Slide_data_12(in_data_to_next_pe_46_12), .Slide_data_13(in_data_to_next_pe_46_13),
                        .Slide_data_14(in_data_to_next_pe_46_14), .Slide_data_15(in_data_to_next_pe_46_15),
                        .Slide_data_16(in_data_to_next_pe_46_16), .Slide_data_17(in_data_to_next_pe_46_17),
                        .Slide_data_18(in_data_to_next_pe_46_18), .Slide_data_19(in_data_to_next_pe_46_19),
                        .Slide_data_20(in_data_to_next_pe_46_20), .Slide_data_21(in_data_to_next_pe_46_21),
                        .Slide_data_22(in_data_to_next_pe_46_22), .Slide_data_23(in_data_to_next_pe_46_23),
                        .Slide_data_24(in_data_to_next_pe_46_24), .Slide_data_25(in_data_to_next_pe_46_25),
                        .Slide_data_26(in_data_to_next_pe_46_26), .Slide_data_27(in_data_to_next_pe_46_27),
                        .Slide_data_28(in_data_to_next_pe_46_28), .Slide_data_29(in_data_to_next_pe_46_29),
                        .Slide_data_30(in_data_to_next_pe_46_30), .Slide_data_31(in_data_to_next_pe_46_31),
                        .result(o_46),
                        .in_data_to_next_pe_0(in_data_to_next_pe_47_0), .in_data_to_next_pe_1(in_data_to_next_pe_47_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_47_2), .in_data_to_next_pe_3(in_data_to_next_pe_47_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_47_4), .in_data_to_next_pe_5(in_data_to_next_pe_47_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_47_6), .in_data_to_next_pe_7(in_data_to_next_pe_47_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_47_8), .in_data_to_next_pe_9(in_data_to_next_pe_47_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_47_10), .in_data_to_next_pe_11(in_data_to_next_pe_47_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_47_12), .in_data_to_next_pe_13(in_data_to_next_pe_47_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_47_14), .in_data_to_next_pe_15(in_data_to_next_pe_47_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_47_16), .in_data_to_next_pe_17(in_data_to_next_pe_47_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_47_18), .in_data_to_next_pe_19(in_data_to_next_pe_47_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_47_20), .in_data_to_next_pe_21(in_data_to_next_pe_47_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_47_22), .in_data_to_next_pe_23(in_data_to_next_pe_47_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_47_24), .in_data_to_next_pe_25(in_data_to_next_pe_47_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_47_26), .in_data_to_next_pe_27(in_data_to_next_pe_47_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_47_28), .in_data_to_next_pe_29(in_data_to_next_pe_47_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_47_30), .in_data_to_next_pe_31(in_data_to_next_pe_47_31),
                        .next_row_en(row_47_en)
        );
        
        PE_Row_B5   PE_R47_B5(   .clk(clk), .rst_n(row_47_en), .new_weight_val(new_weight_val[47]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_47_0), .Slide_data_1(in_data_to_next_pe_47_1),
                        .Slide_data_2(in_data_to_next_pe_47_2), .Slide_data_3(in_data_to_next_pe_47_3),
                        .Slide_data_4(in_data_to_next_pe_47_4), .Slide_data_5(in_data_to_next_pe_47_5),
                        .Slide_data_6(in_data_to_next_pe_47_6), .Slide_data_7(in_data_to_next_pe_47_7),
                        .Slide_data_8(in_data_to_next_pe_47_8), .Slide_data_9(in_data_to_next_pe_47_9),
                        .Slide_data_10(in_data_to_next_pe_47_10), .Slide_data_11(in_data_to_next_pe_47_11),
                        .Slide_data_12(in_data_to_next_pe_47_12), .Slide_data_13(in_data_to_next_pe_47_13),
                        .Slide_data_14(in_data_to_next_pe_47_14), .Slide_data_15(in_data_to_next_pe_47_15),
                        .Slide_data_16(in_data_to_next_pe_47_16), .Slide_data_17(in_data_to_next_pe_47_17),
                        .Slide_data_18(in_data_to_next_pe_47_18), .Slide_data_19(in_data_to_next_pe_47_19),
                        .Slide_data_20(in_data_to_next_pe_47_20), .Slide_data_21(in_data_to_next_pe_47_21),
                        .Slide_data_22(in_data_to_next_pe_47_22), .Slide_data_23(in_data_to_next_pe_47_23),
                        .Slide_data_24(in_data_to_next_pe_47_24), .Slide_data_25(in_data_to_next_pe_47_25),
                        .Slide_data_26(in_data_to_next_pe_47_26), .Slide_data_27(in_data_to_next_pe_47_27),
                        .Slide_data_28(in_data_to_next_pe_47_28), .Slide_data_29(in_data_to_next_pe_47_29),
                        .Slide_data_30(in_data_to_next_pe_47_30), .Slide_data_31(in_data_to_next_pe_47_31),
                        .result(o_47),
                        .in_data_to_next_pe_0(in_data_to_next_pe_48_0), .in_data_to_next_pe_1(in_data_to_next_pe_48_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_48_2), .in_data_to_next_pe_3(in_data_to_next_pe_48_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_48_4), .in_data_to_next_pe_5(in_data_to_next_pe_48_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_48_6), .in_data_to_next_pe_7(in_data_to_next_pe_48_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_48_8), .in_data_to_next_pe_9(in_data_to_next_pe_48_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_48_10), .in_data_to_next_pe_11(in_data_to_next_pe_48_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_48_12), .in_data_to_next_pe_13(in_data_to_next_pe_48_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_48_14), .in_data_to_next_pe_15(in_data_to_next_pe_48_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_48_16), .in_data_to_next_pe_17(in_data_to_next_pe_48_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_48_18), .in_data_to_next_pe_19(in_data_to_next_pe_48_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_48_20), .in_data_to_next_pe_21(in_data_to_next_pe_48_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_48_22), .in_data_to_next_pe_23(in_data_to_next_pe_48_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_48_24), .in_data_to_next_pe_25(in_data_to_next_pe_48_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_48_26), .in_data_to_next_pe_27(in_data_to_next_pe_48_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_48_28), .in_data_to_next_pe_29(in_data_to_next_pe_48_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_48_30), .in_data_to_next_pe_31(in_data_to_next_pe_48_31),
                        .next_row_en(row_48_en)
        );
        
        PE_Row_B5   PE_R48_B5(   .clk(clk), .rst_n(row_48_en), .new_weight_val(new_weight_val[48]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_48_0), .Slide_data_1(in_data_to_next_pe_48_1),
                        .Slide_data_2(in_data_to_next_pe_48_2), .Slide_data_3(in_data_to_next_pe_48_3),
                        .Slide_data_4(in_data_to_next_pe_48_4), .Slide_data_5(in_data_to_next_pe_48_5),
                        .Slide_data_6(in_data_to_next_pe_48_6), .Slide_data_7(in_data_to_next_pe_48_7),
                        .Slide_data_8(in_data_to_next_pe_48_8), .Slide_data_9(in_data_to_next_pe_48_9),
                        .Slide_data_10(in_data_to_next_pe_48_10), .Slide_data_11(in_data_to_next_pe_48_11),
                        .Slide_data_12(in_data_to_next_pe_48_12), .Slide_data_13(in_data_to_next_pe_48_13),
                        .Slide_data_14(in_data_to_next_pe_48_14), .Slide_data_15(in_data_to_next_pe_48_15),
                        .Slide_data_16(in_data_to_next_pe_48_16), .Slide_data_17(in_data_to_next_pe_48_17),
                        .Slide_data_18(in_data_to_next_pe_48_18), .Slide_data_19(in_data_to_next_pe_48_19),
                        .Slide_data_20(in_data_to_next_pe_48_20), .Slide_data_21(in_data_to_next_pe_48_21),
                        .Slide_data_22(in_data_to_next_pe_48_22), .Slide_data_23(in_data_to_next_pe_48_23),
                        .Slide_data_24(in_data_to_next_pe_48_24), .Slide_data_25(in_data_to_next_pe_48_25),
                        .Slide_data_26(in_data_to_next_pe_48_26), .Slide_data_27(in_data_to_next_pe_48_27),
                        .Slide_data_28(in_data_to_next_pe_48_28), .Slide_data_29(in_data_to_next_pe_48_29),
                        .Slide_data_30(in_data_to_next_pe_48_30), .Slide_data_31(in_data_to_next_pe_48_31),
                        .result(o_48),
                        .in_data_to_next_pe_0(in_data_to_next_pe_49_0), .in_data_to_next_pe_1(in_data_to_next_pe_49_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_49_2), .in_data_to_next_pe_3(in_data_to_next_pe_49_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_49_4), .in_data_to_next_pe_5(in_data_to_next_pe_49_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_49_6), .in_data_to_next_pe_7(in_data_to_next_pe_49_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_49_8), .in_data_to_next_pe_9(in_data_to_next_pe_49_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_49_10), .in_data_to_next_pe_11(in_data_to_next_pe_49_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_49_12), .in_data_to_next_pe_13(in_data_to_next_pe_49_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_49_14), .in_data_to_next_pe_15(in_data_to_next_pe_49_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_49_16), .in_data_to_next_pe_17(in_data_to_next_pe_49_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_49_18), .in_data_to_next_pe_19(in_data_to_next_pe_49_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_49_20), .in_data_to_next_pe_21(in_data_to_next_pe_49_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_49_22), .in_data_to_next_pe_23(in_data_to_next_pe_49_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_49_24), .in_data_to_next_pe_25(in_data_to_next_pe_49_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_49_26), .in_data_to_next_pe_27(in_data_to_next_pe_49_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_49_28), .in_data_to_next_pe_29(in_data_to_next_pe_49_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_49_30), .in_data_to_next_pe_31(in_data_to_next_pe_49_31),
                        .next_row_en(row_49_en)
        );
        
        PE_Row_B5   PE_R49_B5(   .clk(clk), .rst_n(row_49_en), .new_weight_val(new_weight_val[49]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_49_0), .Slide_data_1(in_data_to_next_pe_49_1),
                        .Slide_data_2(in_data_to_next_pe_49_2), .Slide_data_3(in_data_to_next_pe_49_3),
                        .Slide_data_4(in_data_to_next_pe_49_4), .Slide_data_5(in_data_to_next_pe_49_5),
                        .Slide_data_6(in_data_to_next_pe_49_6), .Slide_data_7(in_data_to_next_pe_49_7),
                        .Slide_data_8(in_data_to_next_pe_49_8), .Slide_data_9(in_data_to_next_pe_49_9),
                        .Slide_data_10(in_data_to_next_pe_49_10), .Slide_data_11(in_data_to_next_pe_49_11),
                        .Slide_data_12(in_data_to_next_pe_49_12), .Slide_data_13(in_data_to_next_pe_49_13),
                        .Slide_data_14(in_data_to_next_pe_49_14), .Slide_data_15(in_data_to_next_pe_49_15),
                        .Slide_data_16(in_data_to_next_pe_49_16), .Slide_data_17(in_data_to_next_pe_49_17),
                        .Slide_data_18(in_data_to_next_pe_49_18), .Slide_data_19(in_data_to_next_pe_49_19),
                        .Slide_data_20(in_data_to_next_pe_49_20), .Slide_data_21(in_data_to_next_pe_49_21),
                        .Slide_data_22(in_data_to_next_pe_49_22), .Slide_data_23(in_data_to_next_pe_49_23),
                        .Slide_data_24(in_data_to_next_pe_49_24), .Slide_data_25(in_data_to_next_pe_49_25),
                        .Slide_data_26(in_data_to_next_pe_49_26), .Slide_data_27(in_data_to_next_pe_49_27),
                        .Slide_data_28(in_data_to_next_pe_49_28), .Slide_data_29(in_data_to_next_pe_49_29),
                        .Slide_data_30(in_data_to_next_pe_49_30), .Slide_data_31(in_data_to_next_pe_49_31),
                        .result(o_49),
                        .in_data_to_next_pe_0(in_data_to_next_pe_50_0), .in_data_to_next_pe_1(in_data_to_next_pe_50_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_50_2), .in_data_to_next_pe_3(in_data_to_next_pe_50_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_50_4), .in_data_to_next_pe_5(in_data_to_next_pe_50_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_50_6), .in_data_to_next_pe_7(in_data_to_next_pe_50_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_50_8), .in_data_to_next_pe_9(in_data_to_next_pe_50_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_50_10), .in_data_to_next_pe_11(in_data_to_next_pe_50_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_50_12), .in_data_to_next_pe_13(in_data_to_next_pe_50_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_50_14), .in_data_to_next_pe_15(in_data_to_next_pe_50_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_50_16), .in_data_to_next_pe_17(in_data_to_next_pe_50_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_50_18), .in_data_to_next_pe_19(in_data_to_next_pe_50_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_50_20), .in_data_to_next_pe_21(in_data_to_next_pe_50_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_50_22), .in_data_to_next_pe_23(in_data_to_next_pe_50_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_50_24), .in_data_to_next_pe_25(in_data_to_next_pe_50_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_50_26), .in_data_to_next_pe_27(in_data_to_next_pe_50_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_50_28), .in_data_to_next_pe_29(in_data_to_next_pe_50_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_50_30), .in_data_to_next_pe_31(in_data_to_next_pe_50_31),
                        .next_row_en(row_50_en)
        );
        
        PE_Row_B5   PE_R50_B5(   .clk(clk), .rst_n(row_50_en), .new_weight_val(new_weight_val[50]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_50_0), .Slide_data_1(in_data_to_next_pe_50_1),
                        .Slide_data_2(in_data_to_next_pe_50_2), .Slide_data_3(in_data_to_next_pe_50_3),
                        .Slide_data_4(in_data_to_next_pe_50_4), .Slide_data_5(in_data_to_next_pe_50_5),
                        .Slide_data_6(in_data_to_next_pe_50_6), .Slide_data_7(in_data_to_next_pe_50_7),
                        .Slide_data_8(in_data_to_next_pe_50_8), .Slide_data_9(in_data_to_next_pe_50_9),
                        .Slide_data_10(in_data_to_next_pe_50_10), .Slide_data_11(in_data_to_next_pe_50_11),
                        .Slide_data_12(in_data_to_next_pe_50_12), .Slide_data_13(in_data_to_next_pe_50_13),
                        .Slide_data_14(in_data_to_next_pe_50_14), .Slide_data_15(in_data_to_next_pe_50_15),
                        .Slide_data_16(in_data_to_next_pe_50_16), .Slide_data_17(in_data_to_next_pe_50_17),
                        .Slide_data_18(in_data_to_next_pe_50_18), .Slide_data_19(in_data_to_next_pe_50_19),
                        .Slide_data_20(in_data_to_next_pe_50_20), .Slide_data_21(in_data_to_next_pe_50_21),
                        .Slide_data_22(in_data_to_next_pe_50_22), .Slide_data_23(in_data_to_next_pe_50_23),
                        .Slide_data_24(in_data_to_next_pe_50_24), .Slide_data_25(in_data_to_next_pe_50_25),
                        .Slide_data_26(in_data_to_next_pe_50_26), .Slide_data_27(in_data_to_next_pe_50_27),
                        .Slide_data_28(in_data_to_next_pe_50_28), .Slide_data_29(in_data_to_next_pe_50_29),
                        .Slide_data_30(in_data_to_next_pe_50_30), .Slide_data_31(in_data_to_next_pe_50_31),
                        .result(o_50),
                        .in_data_to_next_pe_0(in_data_to_next_pe_51_0), .in_data_to_next_pe_1(in_data_to_next_pe_51_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_51_2), .in_data_to_next_pe_3(in_data_to_next_pe_51_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_51_4), .in_data_to_next_pe_5(in_data_to_next_pe_51_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_51_6), .in_data_to_next_pe_7(in_data_to_next_pe_51_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_51_8), .in_data_to_next_pe_9(in_data_to_next_pe_51_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_51_10), .in_data_to_next_pe_11(in_data_to_next_pe_51_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_51_12), .in_data_to_next_pe_13(in_data_to_next_pe_51_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_51_14), .in_data_to_next_pe_15(in_data_to_next_pe_51_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_51_16), .in_data_to_next_pe_17(in_data_to_next_pe_51_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_51_18), .in_data_to_next_pe_19(in_data_to_next_pe_51_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_51_20), .in_data_to_next_pe_21(in_data_to_next_pe_51_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_51_22), .in_data_to_next_pe_23(in_data_to_next_pe_51_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_51_24), .in_data_to_next_pe_25(in_data_to_next_pe_51_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_51_26), .in_data_to_next_pe_27(in_data_to_next_pe_51_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_51_28), .in_data_to_next_pe_29(in_data_to_next_pe_51_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_51_30), .in_data_to_next_pe_31(in_data_to_next_pe_51_31),
                        .next_row_en(row_51_en)
        );
        
        PE_Row_B5   PE_R51_B5(   .clk(clk), .rst_n(row_51_en), .new_weight_val(new_weight_val[51]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_51_0), .Slide_data_1(in_data_to_next_pe_51_1),
                        .Slide_data_2(in_data_to_next_pe_51_2), .Slide_data_3(in_data_to_next_pe_51_3),
                        .Slide_data_4(in_data_to_next_pe_51_4), .Slide_data_5(in_data_to_next_pe_51_5),
                        .Slide_data_6(in_data_to_next_pe_51_6), .Slide_data_7(in_data_to_next_pe_51_7),
                        .Slide_data_8(in_data_to_next_pe_51_8), .Slide_data_9(in_data_to_next_pe_51_9),
                        .Slide_data_10(in_data_to_next_pe_51_10), .Slide_data_11(in_data_to_next_pe_51_11),
                        .Slide_data_12(in_data_to_next_pe_51_12), .Slide_data_13(in_data_to_next_pe_51_13),
                        .Slide_data_14(in_data_to_next_pe_51_14), .Slide_data_15(in_data_to_next_pe_51_15),
                        .Slide_data_16(in_data_to_next_pe_51_16), .Slide_data_17(in_data_to_next_pe_51_17),
                        .Slide_data_18(in_data_to_next_pe_51_18), .Slide_data_19(in_data_to_next_pe_51_19),
                        .Slide_data_20(in_data_to_next_pe_51_20), .Slide_data_21(in_data_to_next_pe_51_21),
                        .Slide_data_22(in_data_to_next_pe_51_22), .Slide_data_23(in_data_to_next_pe_51_23),
                        .Slide_data_24(in_data_to_next_pe_51_24), .Slide_data_25(in_data_to_next_pe_51_25),
                        .Slide_data_26(in_data_to_next_pe_51_26), .Slide_data_27(in_data_to_next_pe_51_27),
                        .Slide_data_28(in_data_to_next_pe_51_28), .Slide_data_29(in_data_to_next_pe_51_29),
                        .Slide_data_30(in_data_to_next_pe_51_30), .Slide_data_31(in_data_to_next_pe_51_31),
                        .result(o_51),
                        .in_data_to_next_pe_0(in_data_to_next_pe_52_0), .in_data_to_next_pe_1(in_data_to_next_pe_52_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_52_2), .in_data_to_next_pe_3(in_data_to_next_pe_52_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_52_4), .in_data_to_next_pe_5(in_data_to_next_pe_52_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_52_6), .in_data_to_next_pe_7(in_data_to_next_pe_52_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_52_8), .in_data_to_next_pe_9(in_data_to_next_pe_52_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_52_10), .in_data_to_next_pe_11(in_data_to_next_pe_52_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_52_12), .in_data_to_next_pe_13(in_data_to_next_pe_52_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_52_14), .in_data_to_next_pe_15(in_data_to_next_pe_52_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_52_16), .in_data_to_next_pe_17(in_data_to_next_pe_52_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_52_18), .in_data_to_next_pe_19(in_data_to_next_pe_52_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_52_20), .in_data_to_next_pe_21(in_data_to_next_pe_52_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_52_22), .in_data_to_next_pe_23(in_data_to_next_pe_52_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_52_24), .in_data_to_next_pe_25(in_data_to_next_pe_52_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_52_26), .in_data_to_next_pe_27(in_data_to_next_pe_52_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_52_28), .in_data_to_next_pe_29(in_data_to_next_pe_52_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_52_30), .in_data_to_next_pe_31(in_data_to_next_pe_52_31),
                        .next_row_en(row_52_en)
        );
        
        PE_Row_B5   PE_R52_B5(   .clk(clk), .rst_n(row_52_en), .new_weight_val(new_weight_val[52]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_52_0), .Slide_data_1(in_data_to_next_pe_52_1),
                        .Slide_data_2(in_data_to_next_pe_52_2), .Slide_data_3(in_data_to_next_pe_52_3),
                        .Slide_data_4(in_data_to_next_pe_52_4), .Slide_data_5(in_data_to_next_pe_52_5),
                        .Slide_data_6(in_data_to_next_pe_52_6), .Slide_data_7(in_data_to_next_pe_52_7),
                        .Slide_data_8(in_data_to_next_pe_52_8), .Slide_data_9(in_data_to_next_pe_52_9),
                        .Slide_data_10(in_data_to_next_pe_52_10), .Slide_data_11(in_data_to_next_pe_52_11),
                        .Slide_data_12(in_data_to_next_pe_52_12), .Slide_data_13(in_data_to_next_pe_52_13),
                        .Slide_data_14(in_data_to_next_pe_52_14), .Slide_data_15(in_data_to_next_pe_52_15),
                        .Slide_data_16(in_data_to_next_pe_52_16), .Slide_data_17(in_data_to_next_pe_52_17),
                        .Slide_data_18(in_data_to_next_pe_52_18), .Slide_data_19(in_data_to_next_pe_52_19),
                        .Slide_data_20(in_data_to_next_pe_52_20), .Slide_data_21(in_data_to_next_pe_52_21),
                        .Slide_data_22(in_data_to_next_pe_52_22), .Slide_data_23(in_data_to_next_pe_52_23),
                        .Slide_data_24(in_data_to_next_pe_52_24), .Slide_data_25(in_data_to_next_pe_52_25),
                        .Slide_data_26(in_data_to_next_pe_52_26), .Slide_data_27(in_data_to_next_pe_52_27),
                        .Slide_data_28(in_data_to_next_pe_52_28), .Slide_data_29(in_data_to_next_pe_52_29),
                        .Slide_data_30(in_data_to_next_pe_52_30), .Slide_data_31(in_data_to_next_pe_52_31),
                        .result(o_52),
                        .in_data_to_next_pe_0(in_data_to_next_pe_53_0), .in_data_to_next_pe_1(in_data_to_next_pe_53_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_53_2), .in_data_to_next_pe_3(in_data_to_next_pe_53_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_53_4), .in_data_to_next_pe_5(in_data_to_next_pe_53_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_53_6), .in_data_to_next_pe_7(in_data_to_next_pe_53_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_53_8), .in_data_to_next_pe_9(in_data_to_next_pe_53_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_53_10), .in_data_to_next_pe_11(in_data_to_next_pe_53_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_53_12), .in_data_to_next_pe_13(in_data_to_next_pe_53_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_53_14), .in_data_to_next_pe_15(in_data_to_next_pe_53_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_53_16), .in_data_to_next_pe_17(in_data_to_next_pe_53_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_53_18), .in_data_to_next_pe_19(in_data_to_next_pe_53_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_53_20), .in_data_to_next_pe_21(in_data_to_next_pe_53_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_53_22), .in_data_to_next_pe_23(in_data_to_next_pe_53_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_53_24), .in_data_to_next_pe_25(in_data_to_next_pe_53_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_53_26), .in_data_to_next_pe_27(in_data_to_next_pe_53_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_53_28), .in_data_to_next_pe_29(in_data_to_next_pe_53_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_53_30), .in_data_to_next_pe_31(in_data_to_next_pe_53_31),
                        .next_row_en(row_53_en)
        );
        
        PE_Row_B5   PE_R53_B5(   .clk(clk), .rst_n(row_53_en), .new_weight_val(new_weight_val[53]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_53_0), .Slide_data_1(in_data_to_next_pe_53_1),
                        .Slide_data_2(in_data_to_next_pe_53_2), .Slide_data_3(in_data_to_next_pe_53_3),
                        .Slide_data_4(in_data_to_next_pe_53_4), .Slide_data_5(in_data_to_next_pe_53_5),
                        .Slide_data_6(in_data_to_next_pe_53_6), .Slide_data_7(in_data_to_next_pe_53_7),
                        .Slide_data_8(in_data_to_next_pe_53_8), .Slide_data_9(in_data_to_next_pe_53_9),
                        .Slide_data_10(in_data_to_next_pe_53_10), .Slide_data_11(in_data_to_next_pe_53_11),
                        .Slide_data_12(in_data_to_next_pe_53_12), .Slide_data_13(in_data_to_next_pe_53_13),
                        .Slide_data_14(in_data_to_next_pe_53_14), .Slide_data_15(in_data_to_next_pe_53_15),
                        .Slide_data_16(in_data_to_next_pe_53_16), .Slide_data_17(in_data_to_next_pe_53_17),
                        .Slide_data_18(in_data_to_next_pe_53_18), .Slide_data_19(in_data_to_next_pe_53_19),
                        .Slide_data_20(in_data_to_next_pe_53_20), .Slide_data_21(in_data_to_next_pe_53_21),
                        .Slide_data_22(in_data_to_next_pe_53_22), .Slide_data_23(in_data_to_next_pe_53_23),
                        .Slide_data_24(in_data_to_next_pe_53_24), .Slide_data_25(in_data_to_next_pe_53_25),
                        .Slide_data_26(in_data_to_next_pe_53_26), .Slide_data_27(in_data_to_next_pe_53_27),
                        .Slide_data_28(in_data_to_next_pe_53_28), .Slide_data_29(in_data_to_next_pe_53_29),
                        .Slide_data_30(in_data_to_next_pe_53_30), .Slide_data_31(in_data_to_next_pe_53_31),
                        .result(o_53),
                        .in_data_to_next_pe_0(in_data_to_next_pe_54_0), .in_data_to_next_pe_1(in_data_to_next_pe_54_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_54_2), .in_data_to_next_pe_3(in_data_to_next_pe_54_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_54_4), .in_data_to_next_pe_5(in_data_to_next_pe_54_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_54_6), .in_data_to_next_pe_7(in_data_to_next_pe_54_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_54_8), .in_data_to_next_pe_9(in_data_to_next_pe_54_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_54_10), .in_data_to_next_pe_11(in_data_to_next_pe_54_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_54_12), .in_data_to_next_pe_13(in_data_to_next_pe_54_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_54_14), .in_data_to_next_pe_15(in_data_to_next_pe_54_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_54_16), .in_data_to_next_pe_17(in_data_to_next_pe_54_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_54_18), .in_data_to_next_pe_19(in_data_to_next_pe_54_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_54_20), .in_data_to_next_pe_21(in_data_to_next_pe_54_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_54_22), .in_data_to_next_pe_23(in_data_to_next_pe_54_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_54_24), .in_data_to_next_pe_25(in_data_to_next_pe_54_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_54_26), .in_data_to_next_pe_27(in_data_to_next_pe_54_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_54_28), .in_data_to_next_pe_29(in_data_to_next_pe_54_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_54_30), .in_data_to_next_pe_31(in_data_to_next_pe_54_31),
                        .next_row_en(row_54_en)
        );
        
        PE_Row_B5   PE_R54_B5(   .clk(clk), .rst_n(row_54_en), .new_weight_val(new_weight_val[54]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_54_0), .Slide_data_1(in_data_to_next_pe_54_1),
                        .Slide_data_2(in_data_to_next_pe_54_2), .Slide_data_3(in_data_to_next_pe_54_3),
                        .Slide_data_4(in_data_to_next_pe_54_4), .Slide_data_5(in_data_to_next_pe_54_5),
                        .Slide_data_6(in_data_to_next_pe_54_6), .Slide_data_7(in_data_to_next_pe_54_7),
                        .Slide_data_8(in_data_to_next_pe_54_8), .Slide_data_9(in_data_to_next_pe_54_9),
                        .Slide_data_10(in_data_to_next_pe_54_10), .Slide_data_11(in_data_to_next_pe_54_11),
                        .Slide_data_12(in_data_to_next_pe_54_12), .Slide_data_13(in_data_to_next_pe_54_13),
                        .Slide_data_14(in_data_to_next_pe_54_14), .Slide_data_15(in_data_to_next_pe_54_15),
                        .Slide_data_16(in_data_to_next_pe_54_16), .Slide_data_17(in_data_to_next_pe_54_17),
                        .Slide_data_18(in_data_to_next_pe_54_18), .Slide_data_19(in_data_to_next_pe_54_19),
                        .Slide_data_20(in_data_to_next_pe_54_20), .Slide_data_21(in_data_to_next_pe_54_21),
                        .Slide_data_22(in_data_to_next_pe_54_22), .Slide_data_23(in_data_to_next_pe_54_23),
                        .Slide_data_24(in_data_to_next_pe_54_24), .Slide_data_25(in_data_to_next_pe_54_25),
                        .Slide_data_26(in_data_to_next_pe_54_26), .Slide_data_27(in_data_to_next_pe_54_27),
                        .Slide_data_28(in_data_to_next_pe_54_28), .Slide_data_29(in_data_to_next_pe_54_29),
                        .Slide_data_30(in_data_to_next_pe_54_30), .Slide_data_31(in_data_to_next_pe_54_31),
                        .result(o_54),
                        .in_data_to_next_pe_0(in_data_to_next_pe_55_0), .in_data_to_next_pe_1(in_data_to_next_pe_55_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_55_2), .in_data_to_next_pe_3(in_data_to_next_pe_55_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_55_4), .in_data_to_next_pe_5(in_data_to_next_pe_55_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_55_6), .in_data_to_next_pe_7(in_data_to_next_pe_55_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_55_8), .in_data_to_next_pe_9(in_data_to_next_pe_55_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_55_10), .in_data_to_next_pe_11(in_data_to_next_pe_55_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_55_12), .in_data_to_next_pe_13(in_data_to_next_pe_55_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_55_14), .in_data_to_next_pe_15(in_data_to_next_pe_55_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_55_16), .in_data_to_next_pe_17(in_data_to_next_pe_55_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_55_18), .in_data_to_next_pe_19(in_data_to_next_pe_55_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_55_20), .in_data_to_next_pe_21(in_data_to_next_pe_55_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_55_22), .in_data_to_next_pe_23(in_data_to_next_pe_55_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_55_24), .in_data_to_next_pe_25(in_data_to_next_pe_55_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_55_26), .in_data_to_next_pe_27(in_data_to_next_pe_55_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_55_28), .in_data_to_next_pe_29(in_data_to_next_pe_55_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_55_30), .in_data_to_next_pe_31(in_data_to_next_pe_55_31),
                        .next_row_en(row_55_en)
        );
        
        PE_Row_B5   PE_R55_B5(   .clk(clk), .rst_n(row_55_en), .new_weight_val(new_weight_val[55]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_55_0), .Slide_data_1(in_data_to_next_pe_55_1),
                        .Slide_data_2(in_data_to_next_pe_55_2), .Slide_data_3(in_data_to_next_pe_55_3),
                        .Slide_data_4(in_data_to_next_pe_55_4), .Slide_data_5(in_data_to_next_pe_55_5),
                        .Slide_data_6(in_data_to_next_pe_55_6), .Slide_data_7(in_data_to_next_pe_55_7),
                        .Slide_data_8(in_data_to_next_pe_55_8), .Slide_data_9(in_data_to_next_pe_55_9),
                        .Slide_data_10(in_data_to_next_pe_55_10), .Slide_data_11(in_data_to_next_pe_55_11),
                        .Slide_data_12(in_data_to_next_pe_55_12), .Slide_data_13(in_data_to_next_pe_55_13),
                        .Slide_data_14(in_data_to_next_pe_55_14), .Slide_data_15(in_data_to_next_pe_55_15),
                        .Slide_data_16(in_data_to_next_pe_55_16), .Slide_data_17(in_data_to_next_pe_55_17),
                        .Slide_data_18(in_data_to_next_pe_55_18), .Slide_data_19(in_data_to_next_pe_55_19),
                        .Slide_data_20(in_data_to_next_pe_55_20), .Slide_data_21(in_data_to_next_pe_55_21),
                        .Slide_data_22(in_data_to_next_pe_55_22), .Slide_data_23(in_data_to_next_pe_55_23),
                        .Slide_data_24(in_data_to_next_pe_55_24), .Slide_data_25(in_data_to_next_pe_55_25),
                        .Slide_data_26(in_data_to_next_pe_55_26), .Slide_data_27(in_data_to_next_pe_55_27),
                        .Slide_data_28(in_data_to_next_pe_55_28), .Slide_data_29(in_data_to_next_pe_55_29),
                        .Slide_data_30(in_data_to_next_pe_55_30), .Slide_data_31(in_data_to_next_pe_55_31),
                        .result(o_55),
                        .in_data_to_next_pe_0(in_data_to_next_pe_56_0), .in_data_to_next_pe_1(in_data_to_next_pe_56_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_56_2), .in_data_to_next_pe_3(in_data_to_next_pe_56_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_56_4), .in_data_to_next_pe_5(in_data_to_next_pe_56_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_56_6), .in_data_to_next_pe_7(in_data_to_next_pe_56_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_56_8), .in_data_to_next_pe_9(in_data_to_next_pe_56_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_56_10), .in_data_to_next_pe_11(in_data_to_next_pe_56_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_56_12), .in_data_to_next_pe_13(in_data_to_next_pe_56_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_56_14), .in_data_to_next_pe_15(in_data_to_next_pe_56_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_56_16), .in_data_to_next_pe_17(in_data_to_next_pe_56_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_56_18), .in_data_to_next_pe_19(in_data_to_next_pe_56_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_56_20), .in_data_to_next_pe_21(in_data_to_next_pe_56_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_56_22), .in_data_to_next_pe_23(in_data_to_next_pe_56_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_56_24), .in_data_to_next_pe_25(in_data_to_next_pe_56_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_56_26), .in_data_to_next_pe_27(in_data_to_next_pe_56_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_56_28), .in_data_to_next_pe_29(in_data_to_next_pe_56_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_56_30), .in_data_to_next_pe_31(in_data_to_next_pe_56_31),
                        .next_row_en(row_56_en)
        );
        
        PE_Row_B5   PE_R56_B5(   .clk(clk), .rst_n(row_56_en), .new_weight_val(new_weight_val[56]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_56_0), .Slide_data_1(in_data_to_next_pe_56_1),
                        .Slide_data_2(in_data_to_next_pe_56_2), .Slide_data_3(in_data_to_next_pe_56_3),
                        .Slide_data_4(in_data_to_next_pe_56_4), .Slide_data_5(in_data_to_next_pe_56_5),
                        .Slide_data_6(in_data_to_next_pe_56_6), .Slide_data_7(in_data_to_next_pe_56_7),
                        .Slide_data_8(in_data_to_next_pe_56_8), .Slide_data_9(in_data_to_next_pe_56_9),
                        .Slide_data_10(in_data_to_next_pe_56_10), .Slide_data_11(in_data_to_next_pe_56_11),
                        .Slide_data_12(in_data_to_next_pe_56_12), .Slide_data_13(in_data_to_next_pe_56_13),
                        .Slide_data_14(in_data_to_next_pe_56_14), .Slide_data_15(in_data_to_next_pe_56_15),
                        .Slide_data_16(in_data_to_next_pe_56_16), .Slide_data_17(in_data_to_next_pe_56_17),
                        .Slide_data_18(in_data_to_next_pe_56_18), .Slide_data_19(in_data_to_next_pe_56_19),
                        .Slide_data_20(in_data_to_next_pe_56_20), .Slide_data_21(in_data_to_next_pe_56_21),
                        .Slide_data_22(in_data_to_next_pe_56_22), .Slide_data_23(in_data_to_next_pe_56_23),
                        .Slide_data_24(in_data_to_next_pe_56_24), .Slide_data_25(in_data_to_next_pe_56_25),
                        .Slide_data_26(in_data_to_next_pe_56_26), .Slide_data_27(in_data_to_next_pe_56_27),
                        .Slide_data_28(in_data_to_next_pe_56_28), .Slide_data_29(in_data_to_next_pe_56_29),
                        .Slide_data_30(in_data_to_next_pe_56_30), .Slide_data_31(in_data_to_next_pe_56_31),
                        .result(o_56),
                        .in_data_to_next_pe_0(in_data_to_next_pe_57_0), .in_data_to_next_pe_1(in_data_to_next_pe_57_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_57_2), .in_data_to_next_pe_3(in_data_to_next_pe_57_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_57_4), .in_data_to_next_pe_5(in_data_to_next_pe_57_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_57_6), .in_data_to_next_pe_7(in_data_to_next_pe_57_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_57_8), .in_data_to_next_pe_9(in_data_to_next_pe_57_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_57_10), .in_data_to_next_pe_11(in_data_to_next_pe_57_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_57_12), .in_data_to_next_pe_13(in_data_to_next_pe_57_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_57_14), .in_data_to_next_pe_15(in_data_to_next_pe_57_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_57_16), .in_data_to_next_pe_17(in_data_to_next_pe_57_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_57_18), .in_data_to_next_pe_19(in_data_to_next_pe_57_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_57_20), .in_data_to_next_pe_21(in_data_to_next_pe_57_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_57_22), .in_data_to_next_pe_23(in_data_to_next_pe_57_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_57_24), .in_data_to_next_pe_25(in_data_to_next_pe_57_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_57_26), .in_data_to_next_pe_27(in_data_to_next_pe_57_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_57_28), .in_data_to_next_pe_29(in_data_to_next_pe_57_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_57_30), .in_data_to_next_pe_31(in_data_to_next_pe_57_31),
                        .next_row_en(row_57_en)
        );
        
        PE_Row_B5   PE_R57_B5(   .clk(clk), .rst_n(row_57_en), .new_weight_val(new_weight_val[57]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_57_0), .Slide_data_1(in_data_to_next_pe_57_1),
                        .Slide_data_2(in_data_to_next_pe_57_2), .Slide_data_3(in_data_to_next_pe_57_3),
                        .Slide_data_4(in_data_to_next_pe_57_4), .Slide_data_5(in_data_to_next_pe_57_5),
                        .Slide_data_6(in_data_to_next_pe_57_6), .Slide_data_7(in_data_to_next_pe_57_7),
                        .Slide_data_8(in_data_to_next_pe_57_8), .Slide_data_9(in_data_to_next_pe_57_9),
                        .Slide_data_10(in_data_to_next_pe_57_10), .Slide_data_11(in_data_to_next_pe_57_11),
                        .Slide_data_12(in_data_to_next_pe_57_12), .Slide_data_13(in_data_to_next_pe_57_13),
                        .Slide_data_14(in_data_to_next_pe_57_14), .Slide_data_15(in_data_to_next_pe_57_15),
                        .Slide_data_16(in_data_to_next_pe_57_16), .Slide_data_17(in_data_to_next_pe_57_17),
                        .Slide_data_18(in_data_to_next_pe_57_18), .Slide_data_19(in_data_to_next_pe_57_19),
                        .Slide_data_20(in_data_to_next_pe_57_20), .Slide_data_21(in_data_to_next_pe_57_21),
                        .Slide_data_22(in_data_to_next_pe_57_22), .Slide_data_23(in_data_to_next_pe_57_23),
                        .Slide_data_24(in_data_to_next_pe_57_24), .Slide_data_25(in_data_to_next_pe_57_25),
                        .Slide_data_26(in_data_to_next_pe_57_26), .Slide_data_27(in_data_to_next_pe_57_27),
                        .Slide_data_28(in_data_to_next_pe_57_28), .Slide_data_29(in_data_to_next_pe_57_29),
                        .Slide_data_30(in_data_to_next_pe_57_30), .Slide_data_31(in_data_to_next_pe_57_31),
                        .result(o_57),
                        .in_data_to_next_pe_0(in_data_to_next_pe_58_0), .in_data_to_next_pe_1(in_data_to_next_pe_58_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_58_2), .in_data_to_next_pe_3(in_data_to_next_pe_58_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_58_4), .in_data_to_next_pe_5(in_data_to_next_pe_58_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_58_6), .in_data_to_next_pe_7(in_data_to_next_pe_58_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_58_8), .in_data_to_next_pe_9(in_data_to_next_pe_58_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_58_10), .in_data_to_next_pe_11(in_data_to_next_pe_58_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_58_12), .in_data_to_next_pe_13(in_data_to_next_pe_58_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_58_14), .in_data_to_next_pe_15(in_data_to_next_pe_58_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_58_16), .in_data_to_next_pe_17(in_data_to_next_pe_58_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_58_18), .in_data_to_next_pe_19(in_data_to_next_pe_58_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_58_20), .in_data_to_next_pe_21(in_data_to_next_pe_58_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_58_22), .in_data_to_next_pe_23(in_data_to_next_pe_58_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_58_24), .in_data_to_next_pe_25(in_data_to_next_pe_58_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_58_26), .in_data_to_next_pe_27(in_data_to_next_pe_58_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_58_28), .in_data_to_next_pe_29(in_data_to_next_pe_58_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_58_30), .in_data_to_next_pe_31(in_data_to_next_pe_58_31),
                        .next_row_en(row_58_en)
        );
        
        PE_Row_B5   PE_R58_B5(   .clk(clk), .rst_n(row_58_en), .new_weight_val(new_weight_val[58]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_58_0), .Slide_data_1(in_data_to_next_pe_58_1),
                        .Slide_data_2(in_data_to_next_pe_58_2), .Slide_data_3(in_data_to_next_pe_58_3),
                        .Slide_data_4(in_data_to_next_pe_58_4), .Slide_data_5(in_data_to_next_pe_58_5),
                        .Slide_data_6(in_data_to_next_pe_58_6), .Slide_data_7(in_data_to_next_pe_58_7),
                        .Slide_data_8(in_data_to_next_pe_58_8), .Slide_data_9(in_data_to_next_pe_58_9),
                        .Slide_data_10(in_data_to_next_pe_58_10), .Slide_data_11(in_data_to_next_pe_58_11),
                        .Slide_data_12(in_data_to_next_pe_58_12), .Slide_data_13(in_data_to_next_pe_58_13),
                        .Slide_data_14(in_data_to_next_pe_58_14), .Slide_data_15(in_data_to_next_pe_58_15),
                        .Slide_data_16(in_data_to_next_pe_58_16), .Slide_data_17(in_data_to_next_pe_58_17),
                        .Slide_data_18(in_data_to_next_pe_58_18), .Slide_data_19(in_data_to_next_pe_58_19),
                        .Slide_data_20(in_data_to_next_pe_58_20), .Slide_data_21(in_data_to_next_pe_58_21),
                        .Slide_data_22(in_data_to_next_pe_58_22), .Slide_data_23(in_data_to_next_pe_58_23),
                        .Slide_data_24(in_data_to_next_pe_58_24), .Slide_data_25(in_data_to_next_pe_58_25),
                        .Slide_data_26(in_data_to_next_pe_58_26), .Slide_data_27(in_data_to_next_pe_58_27),
                        .Slide_data_28(in_data_to_next_pe_58_28), .Slide_data_29(in_data_to_next_pe_58_29),
                        .Slide_data_30(in_data_to_next_pe_58_30), .Slide_data_31(in_data_to_next_pe_58_31),
                        .result(o_58),
                        .in_data_to_next_pe_0(in_data_to_next_pe_59_0), .in_data_to_next_pe_1(in_data_to_next_pe_59_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_59_2), .in_data_to_next_pe_3(in_data_to_next_pe_59_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_59_4), .in_data_to_next_pe_5(in_data_to_next_pe_59_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_59_6), .in_data_to_next_pe_7(in_data_to_next_pe_59_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_59_8), .in_data_to_next_pe_9(in_data_to_next_pe_59_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_59_10), .in_data_to_next_pe_11(in_data_to_next_pe_59_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_59_12), .in_data_to_next_pe_13(in_data_to_next_pe_59_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_59_14), .in_data_to_next_pe_15(in_data_to_next_pe_59_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_59_16), .in_data_to_next_pe_17(in_data_to_next_pe_59_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_59_18), .in_data_to_next_pe_19(in_data_to_next_pe_59_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_59_20), .in_data_to_next_pe_21(in_data_to_next_pe_59_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_59_22), .in_data_to_next_pe_23(in_data_to_next_pe_59_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_59_24), .in_data_to_next_pe_25(in_data_to_next_pe_59_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_59_26), .in_data_to_next_pe_27(in_data_to_next_pe_59_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_59_28), .in_data_to_next_pe_29(in_data_to_next_pe_59_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_59_30), .in_data_to_next_pe_31(in_data_to_next_pe_59_31),
                        .next_row_en(row_59_en)
        );
        
        PE_Row_B5   PE_R59_B5(   .clk(clk), .rst_n(row_59_en), .new_weight_val(new_weight_val[59]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_59_0), .Slide_data_1(in_data_to_next_pe_59_1),
                        .Slide_data_2(in_data_to_next_pe_59_2), .Slide_data_3(in_data_to_next_pe_59_3),
                        .Slide_data_4(in_data_to_next_pe_59_4), .Slide_data_5(in_data_to_next_pe_59_5),
                        .Slide_data_6(in_data_to_next_pe_59_6), .Slide_data_7(in_data_to_next_pe_59_7),
                        .Slide_data_8(in_data_to_next_pe_59_8), .Slide_data_9(in_data_to_next_pe_59_9),
                        .Slide_data_10(in_data_to_next_pe_59_10), .Slide_data_11(in_data_to_next_pe_59_11),
                        .Slide_data_12(in_data_to_next_pe_59_12), .Slide_data_13(in_data_to_next_pe_59_13),
                        .Slide_data_14(in_data_to_next_pe_59_14), .Slide_data_15(in_data_to_next_pe_59_15),
                        .Slide_data_16(in_data_to_next_pe_59_16), .Slide_data_17(in_data_to_next_pe_59_17),
                        .Slide_data_18(in_data_to_next_pe_59_18), .Slide_data_19(in_data_to_next_pe_59_19),
                        .Slide_data_20(in_data_to_next_pe_59_20), .Slide_data_21(in_data_to_next_pe_59_21),
                        .Slide_data_22(in_data_to_next_pe_59_22), .Slide_data_23(in_data_to_next_pe_59_23),
                        .Slide_data_24(in_data_to_next_pe_59_24), .Slide_data_25(in_data_to_next_pe_59_25),
                        .Slide_data_26(in_data_to_next_pe_59_26), .Slide_data_27(in_data_to_next_pe_59_27),
                        .Slide_data_28(in_data_to_next_pe_59_28), .Slide_data_29(in_data_to_next_pe_59_29),
                        .Slide_data_30(in_data_to_next_pe_59_30), .Slide_data_31(in_data_to_next_pe_59_31),
                        .result(o_59),
                        .in_data_to_next_pe_0(in_data_to_next_pe_60_0), .in_data_to_next_pe_1(in_data_to_next_pe_60_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_60_2), .in_data_to_next_pe_3(in_data_to_next_pe_60_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_60_4), .in_data_to_next_pe_5(in_data_to_next_pe_60_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_60_6), .in_data_to_next_pe_7(in_data_to_next_pe_60_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_60_8), .in_data_to_next_pe_9(in_data_to_next_pe_60_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_60_10), .in_data_to_next_pe_11(in_data_to_next_pe_60_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_60_12), .in_data_to_next_pe_13(in_data_to_next_pe_60_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_60_14), .in_data_to_next_pe_15(in_data_to_next_pe_60_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_60_16), .in_data_to_next_pe_17(in_data_to_next_pe_60_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_60_18), .in_data_to_next_pe_19(in_data_to_next_pe_60_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_60_20), .in_data_to_next_pe_21(in_data_to_next_pe_60_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_60_22), .in_data_to_next_pe_23(in_data_to_next_pe_60_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_60_24), .in_data_to_next_pe_25(in_data_to_next_pe_60_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_60_26), .in_data_to_next_pe_27(in_data_to_next_pe_60_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_60_28), .in_data_to_next_pe_29(in_data_to_next_pe_60_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_60_30), .in_data_to_next_pe_31(in_data_to_next_pe_60_31),
                        .next_row_en(row_60_en)
        );
        
        PE_Row_B5   PE_R60_B5(   .clk(clk), .rst_n(row_60_en), .new_weight_val(new_weight_val[60]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_60_0), .Slide_data_1(in_data_to_next_pe_60_1),
                        .Slide_data_2(in_data_to_next_pe_60_2), .Slide_data_3(in_data_to_next_pe_60_3),
                        .Slide_data_4(in_data_to_next_pe_60_4), .Slide_data_5(in_data_to_next_pe_60_5),
                        .Slide_data_6(in_data_to_next_pe_60_6), .Slide_data_7(in_data_to_next_pe_60_7),
                        .Slide_data_8(in_data_to_next_pe_60_8), .Slide_data_9(in_data_to_next_pe_60_9),
                        .Slide_data_10(in_data_to_next_pe_60_10), .Slide_data_11(in_data_to_next_pe_60_11),
                        .Slide_data_12(in_data_to_next_pe_60_12), .Slide_data_13(in_data_to_next_pe_60_13),
                        .Slide_data_14(in_data_to_next_pe_60_14), .Slide_data_15(in_data_to_next_pe_60_15),
                        .Slide_data_16(in_data_to_next_pe_60_16), .Slide_data_17(in_data_to_next_pe_60_17),
                        .Slide_data_18(in_data_to_next_pe_60_18), .Slide_data_19(in_data_to_next_pe_60_19),
                        .Slide_data_20(in_data_to_next_pe_60_20), .Slide_data_21(in_data_to_next_pe_60_21),
                        .Slide_data_22(in_data_to_next_pe_60_22), .Slide_data_23(in_data_to_next_pe_60_23),
                        .Slide_data_24(in_data_to_next_pe_60_24), .Slide_data_25(in_data_to_next_pe_60_25),
                        .Slide_data_26(in_data_to_next_pe_60_26), .Slide_data_27(in_data_to_next_pe_60_27),
                        .Slide_data_28(in_data_to_next_pe_60_28), .Slide_data_29(in_data_to_next_pe_60_29),
                        .Slide_data_30(in_data_to_next_pe_60_30), .Slide_data_31(in_data_to_next_pe_60_31),
                        .result(o_60),
                        .in_data_to_next_pe_0(in_data_to_next_pe_61_0), .in_data_to_next_pe_1(in_data_to_next_pe_61_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_61_2), .in_data_to_next_pe_3(in_data_to_next_pe_61_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_61_4), .in_data_to_next_pe_5(in_data_to_next_pe_61_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_61_6), .in_data_to_next_pe_7(in_data_to_next_pe_61_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_61_8), .in_data_to_next_pe_9(in_data_to_next_pe_61_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_61_10), .in_data_to_next_pe_11(in_data_to_next_pe_61_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_61_12), .in_data_to_next_pe_13(in_data_to_next_pe_61_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_61_14), .in_data_to_next_pe_15(in_data_to_next_pe_61_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_61_16), .in_data_to_next_pe_17(in_data_to_next_pe_61_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_61_18), .in_data_to_next_pe_19(in_data_to_next_pe_61_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_61_20), .in_data_to_next_pe_21(in_data_to_next_pe_61_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_61_22), .in_data_to_next_pe_23(in_data_to_next_pe_61_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_61_24), .in_data_to_next_pe_25(in_data_to_next_pe_61_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_61_26), .in_data_to_next_pe_27(in_data_to_next_pe_61_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_61_28), .in_data_to_next_pe_29(in_data_to_next_pe_61_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_61_30), .in_data_to_next_pe_31(in_data_to_next_pe_61_31),
                        .next_row_en(row_61_en)
        );
        
        PE_Row_B5   PE_R61_B5(   .clk(clk), .rst_n(row_61_en), .new_weight_val(new_weight_val[61]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_61_0), .Slide_data_1(in_data_to_next_pe_61_1),
                        .Slide_data_2(in_data_to_next_pe_61_2), .Slide_data_3(in_data_to_next_pe_61_3),
                        .Slide_data_4(in_data_to_next_pe_61_4), .Slide_data_5(in_data_to_next_pe_61_5),
                        .Slide_data_6(in_data_to_next_pe_61_6), .Slide_data_7(in_data_to_next_pe_61_7),
                        .Slide_data_8(in_data_to_next_pe_61_8), .Slide_data_9(in_data_to_next_pe_61_9),
                        .Slide_data_10(in_data_to_next_pe_61_10), .Slide_data_11(in_data_to_next_pe_61_11),
                        .Slide_data_12(in_data_to_next_pe_61_12), .Slide_data_13(in_data_to_next_pe_61_13),
                        .Slide_data_14(in_data_to_next_pe_61_14), .Slide_data_15(in_data_to_next_pe_61_15),
                        .Slide_data_16(in_data_to_next_pe_61_16), .Slide_data_17(in_data_to_next_pe_61_17),
                        .Slide_data_18(in_data_to_next_pe_61_18), .Slide_data_19(in_data_to_next_pe_61_19),
                        .Slide_data_20(in_data_to_next_pe_61_20), .Slide_data_21(in_data_to_next_pe_61_21),
                        .Slide_data_22(in_data_to_next_pe_61_22), .Slide_data_23(in_data_to_next_pe_61_23),
                        .Slide_data_24(in_data_to_next_pe_61_24), .Slide_data_25(in_data_to_next_pe_61_25),
                        .Slide_data_26(in_data_to_next_pe_61_26), .Slide_data_27(in_data_to_next_pe_61_27),
                        .Slide_data_28(in_data_to_next_pe_61_28), .Slide_data_29(in_data_to_next_pe_61_29),
                        .Slide_data_30(in_data_to_next_pe_61_30), .Slide_data_31(in_data_to_next_pe_61_31),
                        .result(o_61),
                        .in_data_to_next_pe_0(in_data_to_next_pe_62_0), .in_data_to_next_pe_1(in_data_to_next_pe_62_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_62_2), .in_data_to_next_pe_3(in_data_to_next_pe_62_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_62_4), .in_data_to_next_pe_5(in_data_to_next_pe_62_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_62_6), .in_data_to_next_pe_7(in_data_to_next_pe_62_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_62_8), .in_data_to_next_pe_9(in_data_to_next_pe_62_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_62_10), .in_data_to_next_pe_11(in_data_to_next_pe_62_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_62_12), .in_data_to_next_pe_13(in_data_to_next_pe_62_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_62_14), .in_data_to_next_pe_15(in_data_to_next_pe_62_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_62_16), .in_data_to_next_pe_17(in_data_to_next_pe_62_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_62_18), .in_data_to_next_pe_19(in_data_to_next_pe_62_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_62_20), .in_data_to_next_pe_21(in_data_to_next_pe_62_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_62_22), .in_data_to_next_pe_23(in_data_to_next_pe_62_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_62_24), .in_data_to_next_pe_25(in_data_to_next_pe_62_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_62_26), .in_data_to_next_pe_27(in_data_to_next_pe_62_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_62_28), .in_data_to_next_pe_29(in_data_to_next_pe_62_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_62_30), .in_data_to_next_pe_31(in_data_to_next_pe_62_31),
                        .next_row_en(row_62_en)
        );
        
        PE_Row_B5   PE_R62_B5(   .clk(clk), .rst_n(row_62_en), .new_weight_val(new_weight_val[62]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_62_0), .Slide_data_1(in_data_to_next_pe_62_1),
                        .Slide_data_2(in_data_to_next_pe_62_2), .Slide_data_3(in_data_to_next_pe_62_3),
                        .Slide_data_4(in_data_to_next_pe_62_4), .Slide_data_5(in_data_to_next_pe_62_5),
                        .Slide_data_6(in_data_to_next_pe_62_6), .Slide_data_7(in_data_to_next_pe_62_7),
                        .Slide_data_8(in_data_to_next_pe_62_8), .Slide_data_9(in_data_to_next_pe_62_9),
                        .Slide_data_10(in_data_to_next_pe_62_10), .Slide_data_11(in_data_to_next_pe_62_11),
                        .Slide_data_12(in_data_to_next_pe_62_12), .Slide_data_13(in_data_to_next_pe_62_13),
                        .Slide_data_14(in_data_to_next_pe_62_14), .Slide_data_15(in_data_to_next_pe_62_15),
                        .Slide_data_16(in_data_to_next_pe_62_16), .Slide_data_17(in_data_to_next_pe_62_17),
                        .Slide_data_18(in_data_to_next_pe_62_18), .Slide_data_19(in_data_to_next_pe_62_19),
                        .Slide_data_20(in_data_to_next_pe_62_20), .Slide_data_21(in_data_to_next_pe_62_21),
                        .Slide_data_22(in_data_to_next_pe_62_22), .Slide_data_23(in_data_to_next_pe_62_23),
                        .Slide_data_24(in_data_to_next_pe_62_24), .Slide_data_25(in_data_to_next_pe_62_25),
                        .Slide_data_26(in_data_to_next_pe_62_26), .Slide_data_27(in_data_to_next_pe_62_27),
                        .Slide_data_28(in_data_to_next_pe_62_28), .Slide_data_29(in_data_to_next_pe_62_29),
                        .Slide_data_30(in_data_to_next_pe_62_30), .Slide_data_31(in_data_to_next_pe_62_31),
                        .result(o_62),
                        .in_data_to_next_pe_0(in_data_to_next_pe_63_0), .in_data_to_next_pe_1(in_data_to_next_pe_63_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_63_2), .in_data_to_next_pe_3(in_data_to_next_pe_63_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_63_4), .in_data_to_next_pe_5(in_data_to_next_pe_63_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_63_6), .in_data_to_next_pe_7(in_data_to_next_pe_63_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_63_8), .in_data_to_next_pe_9(in_data_to_next_pe_63_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_63_10), .in_data_to_next_pe_11(in_data_to_next_pe_63_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_63_12), .in_data_to_next_pe_13(in_data_to_next_pe_63_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_63_14), .in_data_to_next_pe_15(in_data_to_next_pe_63_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_63_16), .in_data_to_next_pe_17(in_data_to_next_pe_63_17),
                        .in_data_to_next_pe_18(in_data_to_next_pe_63_18), .in_data_to_next_pe_19(in_data_to_next_pe_63_19),
                        .in_data_to_next_pe_20(in_data_to_next_pe_63_20), .in_data_to_next_pe_21(in_data_to_next_pe_63_21),
                        .in_data_to_next_pe_22(in_data_to_next_pe_63_22), .in_data_to_next_pe_23(in_data_to_next_pe_63_23),
                        .in_data_to_next_pe_24(in_data_to_next_pe_63_24), .in_data_to_next_pe_25(in_data_to_next_pe_63_25),
                        .in_data_to_next_pe_26(in_data_to_next_pe_63_26), .in_data_to_next_pe_27(in_data_to_next_pe_63_27),
                        .in_data_to_next_pe_28(in_data_to_next_pe_63_28), .in_data_to_next_pe_29(in_data_to_next_pe_63_29),
                        .in_data_to_next_pe_30(in_data_to_next_pe_63_30), .in_data_to_next_pe_31(in_data_to_next_pe_63_31),
                        .next_row_en(row_63_en)
        );
        
        PE_Row_B5   PE_R63_B5(   .clk(clk), .rst_n(row_63_en), .new_weight_val(new_weight_val[63]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3),
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11),
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19),
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23),
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27),
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .Slide_data_0(in_data_to_next_pe_63_0), .Slide_data_1(in_data_to_next_pe_63_1),
                        .Slide_data_2(in_data_to_next_pe_63_2), .Slide_data_3(in_data_to_next_pe_63_3),
                        .Slide_data_4(in_data_to_next_pe_63_4), .Slide_data_5(in_data_to_next_pe_63_5),
                        .Slide_data_6(in_data_to_next_pe_63_6), .Slide_data_7(in_data_to_next_pe_63_7),
                        .Slide_data_8(in_data_to_next_pe_63_8), .Slide_data_9(in_data_to_next_pe_63_9),
                        .Slide_data_10(in_data_to_next_pe_63_10), .Slide_data_11(in_data_to_next_pe_63_11),
                        .Slide_data_12(in_data_to_next_pe_63_12), .Slide_data_13(in_data_to_next_pe_63_13),
                        .Slide_data_14(in_data_to_next_pe_63_14), .Slide_data_15(in_data_to_next_pe_63_15),
                        .Slide_data_16(in_data_to_next_pe_63_16), .Slide_data_17(in_data_to_next_pe_63_17),
                        .Slide_data_18(in_data_to_next_pe_63_18), .Slide_data_19(in_data_to_next_pe_63_19),
                        .Slide_data_20(in_data_to_next_pe_63_20), .Slide_data_21(in_data_to_next_pe_63_21),
                        .Slide_data_22(in_data_to_next_pe_63_22), .Slide_data_23(in_data_to_next_pe_63_23),
                        .Slide_data_24(in_data_to_next_pe_63_24), .Slide_data_25(in_data_to_next_pe_63_25),
                        .Slide_data_26(in_data_to_next_pe_63_26), .Slide_data_27(in_data_to_next_pe_63_27),
                        .Slide_data_28(in_data_to_next_pe_63_28), .Slide_data_29(in_data_to_next_pe_63_29),
                        .Slide_data_30(in_data_to_next_pe_63_30), .Slide_data_31(in_data_to_next_pe_63_31),
                        .result(o_63),
                        .in_data_to_next_pe_0(), .in_data_to_next_pe_1(),
                        .in_data_to_next_pe_2(), .in_data_to_next_pe_3(),
                        .in_data_to_next_pe_4(), .in_data_to_next_pe_5(),
                        .in_data_to_next_pe_6(), .in_data_to_next_pe_7(),
                        .in_data_to_next_pe_8(), .in_data_to_next_pe_9(),
                        .in_data_to_next_pe_10(), .in_data_to_next_pe_11(),
                        .in_data_to_next_pe_12(), .in_data_to_next_pe_13(),
                        .in_data_to_next_pe_14(), .in_data_to_next_pe_15(),
                        .in_data_to_next_pe_16(), .in_data_to_next_pe_17(),
                        .in_data_to_next_pe_18(), .in_data_to_next_pe_19(),
                        .in_data_to_next_pe_20(), .in_data_to_next_pe_21(),
                        .in_data_to_next_pe_22(), .in_data_to_next_pe_23(),
                        .in_data_to_next_pe_24(), .in_data_to_next_pe_25(),
                        .in_data_to_next_pe_26(), .in_data_to_next_pe_27(),
                        .in_data_to_next_pe_28(), .in_data_to_next_pe_29(),
                        .in_data_to_next_pe_30(), .in_data_to_next_pe_31(),
                        .next_row_en()
        );
        
        

endmodule
