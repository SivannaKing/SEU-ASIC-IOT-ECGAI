`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/05/08 20:05:52
// Design Name: 
// Module Name: PE_Array_B6
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module PE_Array_B6(
    input                       clk,
    input                       rst_n,
    input               [4:0]   new_weight_val,
    input               [6:0]   w_0, w_1, w_2, w_3, w_4, w_5, w_6, w_7, w_8, w_9, w_10, w_11, w_12, w_13, w_14, w_15,
                                w_16, w_17, w_18, w_19, w_20, w_21, w_22, w_23, w_24, w_25, w_26, w_27, w_28, w_29, w_30, w_31,
                                w_32, w_33, w_34, w_35, w_36, w_37, w_38, w_39, w_40, w_41, w_42, w_43, w_44, w_45, w_46, w_47, 
                                w_48, w_49, w_50, w_51, w_52, w_53, w_54, w_55, w_56, w_57, w_58, w_59, w_60, w_61, w_62, w_63,
    input   wire        [6:0]   Slide_data_0, Slide_data_1, Slide_data_2, Slide_data_3, Slide_data_4, Slide_data_5, Slide_data_6, Slide_data_7,
                                Slide_data_8, Slide_data_9, Slide_data_10, Slide_data_11, Slide_data_12, Slide_data_13, Slide_data_14, Slide_data_15,
                                Slide_data_16, Slide_data_17, Slide_data_18, Slide_data_19, Slide_data_20, Slide_data_21, Slide_data_22, Slide_data_23, 
                                Slide_data_24, Slide_data_25, Slide_data_26, Slide_data_27, Slide_data_28, Slide_data_29, Slide_data_30, Slide_data_31,
                                Slide_data_32, Slide_data_33, Slide_data_34, Slide_data_35, Slide_data_36, Slide_data_37, Slide_data_38, Slide_data_39, 
                                Slide_data_40, Slide_data_41, Slide_data_42, Slide_data_43, Slide_data_44, Slide_data_45, Slide_data_46, Slide_data_47, 
                                Slide_data_48, Slide_data_49, Slide_data_50, Slide_data_51, Slide_data_52, Slide_data_53, Slide_data_54, Slide_data_55, 
                                Slide_data_56, Slide_data_57, Slide_data_58, Slide_data_59, Slide_data_60, Slide_data_61, Slide_data_62, Slide_data_63,
    output  wire signed [9:0]   o_0, o_1, o_2, o_3, o_4,
    output  wire                o_0_val
    );
wire    [6:0]           in_data_to_next_pe_1_0, in_data_to_next_pe_1_1, in_data_to_next_pe_1_2, in_data_to_next_pe_1_3,
                        in_data_to_next_pe_1_4, in_data_to_next_pe_1_5, in_data_to_next_pe_1_6, in_data_to_next_pe_1_7,
                        in_data_to_next_pe_1_8, in_data_to_next_pe_1_9, in_data_to_next_pe_1_10, in_data_to_next_pe_1_11,
                        in_data_to_next_pe_1_12, in_data_to_next_pe_1_13, in_data_to_next_pe_1_14, in_data_to_next_pe_1_15,
                        in_data_to_next_pe_1_16, in_data_to_next_pe_1_17, in_data_to_next_pe_1_18, in_data_to_next_pe_1_19,
                        in_data_to_next_pe_1_20, in_data_to_next_pe_1_21, in_data_to_next_pe_1_22, in_data_to_next_pe_1_23,
                        in_data_to_next_pe_1_24, in_data_to_next_pe_1_25, in_data_to_next_pe_1_26, in_data_to_next_pe_1_27,
                        in_data_to_next_pe_1_28, in_data_to_next_pe_1_29, in_data_to_next_pe_1_30, in_data_to_next_pe_1_31,
                        in_data_to_next_pe_1_32, in_data_to_next_pe_1_33, in_data_to_next_pe_1_34, in_data_to_next_pe_1_35,
                        in_data_to_next_pe_1_36, in_data_to_next_pe_1_37, in_data_to_next_pe_1_38, in_data_to_next_pe_1_39,
                        in_data_to_next_pe_1_40, in_data_to_next_pe_1_41, in_data_to_next_pe_1_42, in_data_to_next_pe_1_43,
                        in_data_to_next_pe_1_44, in_data_to_next_pe_1_45, in_data_to_next_pe_1_46, in_data_to_next_pe_1_47,
                        in_data_to_next_pe_1_48, in_data_to_next_pe_1_49, in_data_to_next_pe_1_50, in_data_to_next_pe_1_51,
                        in_data_to_next_pe_1_52, in_data_to_next_pe_1_53, in_data_to_next_pe_1_54, in_data_to_next_pe_1_55,
                        in_data_to_next_pe_1_56, in_data_to_next_pe_1_57, in_data_to_next_pe_1_58, in_data_to_next_pe_1_59,
                        in_data_to_next_pe_1_60, in_data_to_next_pe_1_61, in_data_to_next_pe_1_62, in_data_to_next_pe_1_63,
                        
                        in_data_to_next_pe_2_0, in_data_to_next_pe_2_1, in_data_to_next_pe_2_2, in_data_to_next_pe_2_3,
                        in_data_to_next_pe_2_4, in_data_to_next_pe_2_5, in_data_to_next_pe_2_6, in_data_to_next_pe_2_7,
                        in_data_to_next_pe_2_8, in_data_to_next_pe_2_9, in_data_to_next_pe_2_10, in_data_to_next_pe_2_11,
                        in_data_to_next_pe_2_12, in_data_to_next_pe_2_13, in_data_to_next_pe_2_14, in_data_to_next_pe_2_15,
                        in_data_to_next_pe_2_16, in_data_to_next_pe_2_17, in_data_to_next_pe_2_18, in_data_to_next_pe_2_19,
                        in_data_to_next_pe_2_20, in_data_to_next_pe_2_21, in_data_to_next_pe_2_22, in_data_to_next_pe_2_23,
                        in_data_to_next_pe_2_24, in_data_to_next_pe_2_25, in_data_to_next_pe_2_26, in_data_to_next_pe_2_27,
                        in_data_to_next_pe_2_28, in_data_to_next_pe_2_29, in_data_to_next_pe_2_30, in_data_to_next_pe_2_31,
                        in_data_to_next_pe_2_32, in_data_to_next_pe_2_33, in_data_to_next_pe_2_34, in_data_to_next_pe_2_35,
                        in_data_to_next_pe_2_36, in_data_to_next_pe_2_37, in_data_to_next_pe_2_38, in_data_to_next_pe_2_39,
                        in_data_to_next_pe_2_40, in_data_to_next_pe_2_41, in_data_to_next_pe_2_42, in_data_to_next_pe_2_43,
                        in_data_to_next_pe_2_44, in_data_to_next_pe_2_45, in_data_to_next_pe_2_46, in_data_to_next_pe_2_47,
                        in_data_to_next_pe_2_48, in_data_to_next_pe_2_49, in_data_to_next_pe_2_50, in_data_to_next_pe_2_51,
                        in_data_to_next_pe_2_52, in_data_to_next_pe_2_53, in_data_to_next_pe_2_54, in_data_to_next_pe_2_55,
                        in_data_to_next_pe_2_56, in_data_to_next_pe_2_57, in_data_to_next_pe_2_58, in_data_to_next_pe_2_59,
                        in_data_to_next_pe_2_60, in_data_to_next_pe_2_61, in_data_to_next_pe_2_62, in_data_to_next_pe_2_63,
                        
                        in_data_to_next_pe_3_0, in_data_to_next_pe_3_1, in_data_to_next_pe_3_2, in_data_to_next_pe_3_3,
                        in_data_to_next_pe_3_4, in_data_to_next_pe_3_5, in_data_to_next_pe_3_6, in_data_to_next_pe_3_7,
                        in_data_to_next_pe_3_8, in_data_to_next_pe_3_9, in_data_to_next_pe_3_10, in_data_to_next_pe_3_11,
                        in_data_to_next_pe_3_12, in_data_to_next_pe_3_13, in_data_to_next_pe_3_14, in_data_to_next_pe_3_15,
                        in_data_to_next_pe_3_16, in_data_to_next_pe_3_17, in_data_to_next_pe_3_18, in_data_to_next_pe_3_19,
                        in_data_to_next_pe_3_20, in_data_to_next_pe_3_21, in_data_to_next_pe_3_22, in_data_to_next_pe_3_23,
                        in_data_to_next_pe_3_24, in_data_to_next_pe_3_25, in_data_to_next_pe_3_26, in_data_to_next_pe_3_27,
                        in_data_to_next_pe_3_28, in_data_to_next_pe_3_29, in_data_to_next_pe_3_30, in_data_to_next_pe_3_31,
                        in_data_to_next_pe_3_32, in_data_to_next_pe_3_33, in_data_to_next_pe_3_34, in_data_to_next_pe_3_35,
                        in_data_to_next_pe_3_36, in_data_to_next_pe_3_37, in_data_to_next_pe_3_38, in_data_to_next_pe_3_39,
                        in_data_to_next_pe_3_40, in_data_to_next_pe_3_41, in_data_to_next_pe_3_42, in_data_to_next_pe_3_43,
                        in_data_to_next_pe_3_44, in_data_to_next_pe_3_45, in_data_to_next_pe_3_46, in_data_to_next_pe_3_47,
                        in_data_to_next_pe_3_48, in_data_to_next_pe_3_49, in_data_to_next_pe_3_50, in_data_to_next_pe_3_51,
                        in_data_to_next_pe_3_52, in_data_to_next_pe_3_53, in_data_to_next_pe_3_54, in_data_to_next_pe_3_55,
                        in_data_to_next_pe_3_56, in_data_to_next_pe_3_57, in_data_to_next_pe_3_58, in_data_to_next_pe_3_59,
                        in_data_to_next_pe_3_60, in_data_to_next_pe_3_61, in_data_to_next_pe_3_62, in_data_to_next_pe_3_63,
                        
                        in_data_to_next_pe_4_0, in_data_to_next_pe_4_1, in_data_to_next_pe_4_2, in_data_to_next_pe_4_3,
                        in_data_to_next_pe_4_4, in_data_to_next_pe_4_5, in_data_to_next_pe_4_6, in_data_to_next_pe_4_7,
                        in_data_to_next_pe_4_8, in_data_to_next_pe_4_9, in_data_to_next_pe_4_10, in_data_to_next_pe_4_11,
                        in_data_to_next_pe_4_12, in_data_to_next_pe_4_13, in_data_to_next_pe_4_14, in_data_to_next_pe_4_15,
                        in_data_to_next_pe_4_16, in_data_to_next_pe_4_17, in_data_to_next_pe_4_18, in_data_to_next_pe_4_19,
                        in_data_to_next_pe_4_20, in_data_to_next_pe_4_21, in_data_to_next_pe_4_22, in_data_to_next_pe_4_23,
                        in_data_to_next_pe_4_24, in_data_to_next_pe_4_25, in_data_to_next_pe_4_26, in_data_to_next_pe_4_27,
                        in_data_to_next_pe_4_28, in_data_to_next_pe_4_29, in_data_to_next_pe_4_30, in_data_to_next_pe_4_31,
                        in_data_to_next_pe_4_32, in_data_to_next_pe_4_33, in_data_to_next_pe_4_34, in_data_to_next_pe_4_35,
                        in_data_to_next_pe_4_36, in_data_to_next_pe_4_37, in_data_to_next_pe_4_38, in_data_to_next_pe_4_39,
                        in_data_to_next_pe_4_40, in_data_to_next_pe_4_41, in_data_to_next_pe_4_42, in_data_to_next_pe_4_43,
                        in_data_to_next_pe_4_44, in_data_to_next_pe_4_45, in_data_to_next_pe_4_46, in_data_to_next_pe_4_47,
                        in_data_to_next_pe_4_48, in_data_to_next_pe_4_49, in_data_to_next_pe_4_50, in_data_to_next_pe_4_51,
                        in_data_to_next_pe_4_52, in_data_to_next_pe_4_53, in_data_to_next_pe_4_54, in_data_to_next_pe_4_55,
                        in_data_to_next_pe_4_56, in_data_to_next_pe_4_57, in_data_to_next_pe_4_58, in_data_to_next_pe_4_59,
                        in_data_to_next_pe_4_60, in_data_to_next_pe_4_61, in_data_to_next_pe_4_62, in_data_to_next_pe_4_63;
wire                    row_1_en, row_2_en,  row_3_en,  row_4_en;        

PE_Row_B6   PE_R0_B6(   .clk(clk), .rst_n(rst_n), .new_weight_val(new_weight_val[0]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3), 
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11), 
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19), 
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23), 
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27), 
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .w_32(w_32), .w_33(w_33), .w_34(w_34), .w_35(w_35), 
                        .w_36(w_36), .w_37(w_37), .w_38(w_38), .w_39(w_39), 
                        .w_40(w_40), .w_41(w_41), .w_42(w_42), .w_43(w_43), 
                        .w_44(w_44), .w_45(w_45), .w_46(w_46), .w_47(w_47), 
                        .w_48(w_48), .w_49(w_49), .w_50(w_50), .w_51(w_51), 
                        .w_52(w_52), .w_53(w_53), .w_54(w_54), .w_55(w_55), 
                        .w_56(w_56), .w_57(w_57), .w_58(w_58), .w_59(w_59), 
                        .w_60(w_60), .w_61(w_61), .w_62(w_62), .w_63(w_63), 
                        .Slide_data_0(Slide_data_0), .Slide_data_1(Slide_data_1),
                        .Slide_data_2(Slide_data_2), .Slide_data_3(Slide_data_3), 
                        .Slide_data_4(Slide_data_4), .Slide_data_5(Slide_data_5),
                        .Slide_data_6(Slide_data_6), .Slide_data_7(Slide_data_7),
                        .Slide_data_8(Slide_data_8), .Slide_data_9(Slide_data_9),
                        .Slide_data_10(Slide_data_10), .Slide_data_11(Slide_data_11), 
                        .Slide_data_12(Slide_data_12), .Slide_data_13(Slide_data_13),
                        .Slide_data_14(Slide_data_14), .Slide_data_15(Slide_data_15),
                        .Slide_data_16(Slide_data_16), .Slide_data_17(Slide_data_17), 
                        .Slide_data_18(Slide_data_18), .Slide_data_19(Slide_data_19), 
                        .Slide_data_20(Slide_data_20), .Slide_data_21(Slide_data_21), 
                        .Slide_data_22(Slide_data_22), .Slide_data_23(Slide_data_23), 
                        .Slide_data_24(Slide_data_24), .Slide_data_25(Slide_data_25), 
                        .Slide_data_26(Slide_data_26), .Slide_data_27(Slide_data_27), 
                        .Slide_data_28(Slide_data_28), .Slide_data_29(Slide_data_29), 
                        .Slide_data_30(Slide_data_30), .Slide_data_31(Slide_data_31), 
                        .Slide_data_32(Slide_data_32), .Slide_data_33(Slide_data_33), 
                        .Slide_data_34(Slide_data_34), .Slide_data_35(Slide_data_35), 
                        .Slide_data_36(Slide_data_36), .Slide_data_37(Slide_data_37), 
                        .Slide_data_38(Slide_data_38), .Slide_data_39(Slide_data_39), 
                        .Slide_data_40(Slide_data_40), .Slide_data_41(Slide_data_41), 
                        .Slide_data_42(Slide_data_42), .Slide_data_43(Slide_data_43), 
                        .Slide_data_44(Slide_data_44), .Slide_data_45(Slide_data_45), 
                        .Slide_data_46(Slide_data_46), .Slide_data_47(Slide_data_47), 
                        .Slide_data_48(Slide_data_48), .Slide_data_49(Slide_data_49), 
                        .Slide_data_50(Slide_data_50), .Slide_data_51(Slide_data_51), 
                        .Slide_data_52(Slide_data_52), .Slide_data_53(Slide_data_53), 
                        .Slide_data_54(Slide_data_54), .Slide_data_55(Slide_data_55), 
                        .Slide_data_56(Slide_data_56), .Slide_data_57(Slide_data_57), 
                        .Slide_data_58(Slide_data_58), .Slide_data_59(Slide_data_59), 
                        .Slide_data_60(Slide_data_60), .Slide_data_61(Slide_data_61), 
                        .Slide_data_62(Slide_data_62), .Slide_data_63(Slide_data_63),
                        .result(o_0),
                        .in_data_to_next_pe_0(in_data_to_next_pe_1_0), .in_data_to_next_pe_1(in_data_to_next_pe_1_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_1_2), .in_data_to_next_pe_3(in_data_to_next_pe_1_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_1_4), .in_data_to_next_pe_5(in_data_to_next_pe_1_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_1_6), .in_data_to_next_pe_7(in_data_to_next_pe_1_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_1_8), .in_data_to_next_pe_9(in_data_to_next_pe_1_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_1_10), .in_data_to_next_pe_11(in_data_to_next_pe_1_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_1_12), .in_data_to_next_pe_13(in_data_to_next_pe_1_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_1_14), .in_data_to_next_pe_15(in_data_to_next_pe_1_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_1_16), .in_data_to_next_pe_17(in_data_to_next_pe_1_17), 
                        .in_data_to_next_pe_18(in_data_to_next_pe_1_18), .in_data_to_next_pe_19(in_data_to_next_pe_1_19), 
                        .in_data_to_next_pe_20(in_data_to_next_pe_1_20), .in_data_to_next_pe_21(in_data_to_next_pe_1_21), 
                        .in_data_to_next_pe_22(in_data_to_next_pe_1_22), .in_data_to_next_pe_23(in_data_to_next_pe_1_23), 
                        .in_data_to_next_pe_24(in_data_to_next_pe_1_24), .in_data_to_next_pe_25(in_data_to_next_pe_1_25), 
                        .in_data_to_next_pe_26(in_data_to_next_pe_1_26), .in_data_to_next_pe_27(in_data_to_next_pe_1_27), 
                        .in_data_to_next_pe_28(in_data_to_next_pe_1_28), .in_data_to_next_pe_29(in_data_to_next_pe_1_29), 
                        .in_data_to_next_pe_30(in_data_to_next_pe_1_30), .in_data_to_next_pe_31(in_data_to_next_pe_1_31),
                        .in_data_to_next_pe_32(in_data_to_next_pe_1_32), .in_data_to_next_pe_33(in_data_to_next_pe_1_33), 
                        .in_data_to_next_pe_34(in_data_to_next_pe_1_34), .in_data_to_next_pe_35(in_data_to_next_pe_1_35), 
                        .in_data_to_next_pe_36(in_data_to_next_pe_1_36), .in_data_to_next_pe_37(in_data_to_next_pe_1_37), 
                        .in_data_to_next_pe_38(in_data_to_next_pe_1_38), .in_data_to_next_pe_39(in_data_to_next_pe_1_39), 
                        .in_data_to_next_pe_40(in_data_to_next_pe_1_40), .in_data_to_next_pe_41(in_data_to_next_pe_1_41), 
                        .in_data_to_next_pe_42(in_data_to_next_pe_1_42), .in_data_to_next_pe_43(in_data_to_next_pe_1_43), 
                        .in_data_to_next_pe_44(in_data_to_next_pe_1_44), .in_data_to_next_pe_45(in_data_to_next_pe_1_45), 
                        .in_data_to_next_pe_46(in_data_to_next_pe_1_46), .in_data_to_next_pe_47(in_data_to_next_pe_1_47), 
                        .in_data_to_next_pe_48(in_data_to_next_pe_1_48), .in_data_to_next_pe_49(in_data_to_next_pe_1_49), 
                        .in_data_to_next_pe_50(in_data_to_next_pe_1_50), .in_data_to_next_pe_51(in_data_to_next_pe_1_51), 
                        .in_data_to_next_pe_52(in_data_to_next_pe_1_52), .in_data_to_next_pe_53(in_data_to_next_pe_1_53), 
                        .in_data_to_next_pe_54(in_data_to_next_pe_1_54), .in_data_to_next_pe_55(in_data_to_next_pe_1_55), 
                        .in_data_to_next_pe_56(in_data_to_next_pe_1_56), .in_data_to_next_pe_57(in_data_to_next_pe_1_57), 
                        .in_data_to_next_pe_58(in_data_to_next_pe_1_58), .in_data_to_next_pe_59(in_data_to_next_pe_1_59), 
                        .in_data_to_next_pe_60(in_data_to_next_pe_1_60), .in_data_to_next_pe_61(in_data_to_next_pe_1_61), 
                        .in_data_to_next_pe_62(in_data_to_next_pe_1_62), .in_data_to_next_pe_63(in_data_to_next_pe_1_63), 
                        .next_row_en(row_1_en),  
                        .out_val(o_0_val)
);      


PE_Row_B6   PE_R1_B6(   .clk(clk), .rst_n(rst_n), .new_weight_val(new_weight_val[1]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3), 
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11), 
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19), 
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23), 
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27), 
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .w_32(w_32), .w_33(w_33), .w_34(w_34), .w_35(w_35), 
                        .w_36(w_36), .w_37(w_37), .w_38(w_38), .w_39(w_39), 
                        .w_40(w_40), .w_41(w_41), .w_42(w_42), .w_43(w_43), 
                        .w_44(w_44), .w_45(w_45), .w_46(w_46), .w_47(w_47), 
                        .w_48(w_48), .w_49(w_49), .w_50(w_50), .w_51(w_51), 
                        .w_52(w_52), .w_53(w_53), .w_54(w_54), .w_55(w_55), 
                        .w_56(w_56), .w_57(w_57), .w_58(w_58), .w_59(w_59), 
                        .w_60(w_60), .w_61(w_61), .w_62(w_62), .w_63(w_63),  
                        .Slide_data_0(in_data_to_next_pe_1_0), .Slide_data_1(in_data_to_next_pe_1_1),
                        .Slide_data_2(in_data_to_next_pe_1_2),.Slide_data_3(in_data_to_next_pe_1_3),
                        .Slide_data_4(in_data_to_next_pe_1_4),.Slide_data_5(in_data_to_next_pe_1_5),
                        .Slide_data_6(in_data_to_next_pe_1_6),.Slide_data_7(in_data_to_next_pe_1_7),
                        .Slide_data_8(in_data_to_next_pe_1_8),.Slide_data_9(in_data_to_next_pe_1_9),
                        .Slide_data_10(in_data_to_next_pe_1_10),.Slide_data_11(in_data_to_next_pe_1_11),
                        .Slide_data_12(in_data_to_next_pe_1_12),.Slide_data_13(in_data_to_next_pe_1_13),
                        .Slide_data_14(in_data_to_next_pe_1_14),.Slide_data_15(in_data_to_next_pe_1_15),
                        .Slide_data_16(in_data_to_next_pe_1_16),.Slide_data_17(in_data_to_next_pe_1_17),
                        .Slide_data_18(in_data_to_next_pe_1_18),.Slide_data_19(in_data_to_next_pe_1_19),
                        .Slide_data_20(in_data_to_next_pe_1_20),.Slide_data_21(in_data_to_next_pe_1_21),
                        .Slide_data_22(in_data_to_next_pe_1_22),.Slide_data_23(in_data_to_next_pe_1_23),
                        .Slide_data_24(in_data_to_next_pe_1_24),.Slide_data_25(in_data_to_next_pe_1_25),
                        .Slide_data_26(in_data_to_next_pe_1_26),.Slide_data_27(in_data_to_next_pe_1_27),
                        .Slide_data_28(in_data_to_next_pe_1_28),.Slide_data_29(in_data_to_next_pe_1_29),
                        .Slide_data_30(in_data_to_next_pe_1_30),.Slide_data_31(in_data_to_next_pe_1_31),
                        .Slide_data_32(in_data_to_next_pe_1_32),.Slide_data_33(in_data_to_next_pe_1_33),
                        .Slide_data_34(in_data_to_next_pe_1_34),.Slide_data_35(in_data_to_next_pe_1_35),
                        .Slide_data_36(in_data_to_next_pe_1_36),.Slide_data_37(in_data_to_next_pe_1_37),
                        .Slide_data_38(in_data_to_next_pe_1_38),.Slide_data_39(in_data_to_next_pe_1_39),
                        .Slide_data_40(in_data_to_next_pe_1_40),.Slide_data_41(in_data_to_next_pe_1_41),
                        .Slide_data_42(in_data_to_next_pe_1_42),.Slide_data_43(in_data_to_next_pe_1_43),
                        .Slide_data_44(in_data_to_next_pe_1_44),.Slide_data_45(in_data_to_next_pe_1_45),
                        .Slide_data_46(in_data_to_next_pe_1_46),.Slide_data_47(in_data_to_next_pe_1_47),
                        .Slide_data_48(in_data_to_next_pe_1_48),.Slide_data_49(in_data_to_next_pe_1_49),
                        .Slide_data_50(in_data_to_next_pe_1_50),.Slide_data_51(in_data_to_next_pe_1_51),
                        .Slide_data_52(in_data_to_next_pe_1_52),.Slide_data_53(in_data_to_next_pe_1_53),
                        .Slide_data_54(in_data_to_next_pe_1_54),.Slide_data_55(in_data_to_next_pe_1_55),
                        .Slide_data_56(in_data_to_next_pe_1_56),.Slide_data_57(in_data_to_next_pe_1_57),
                        .Slide_data_58(in_data_to_next_pe_1_58),.Slide_data_59(in_data_to_next_pe_1_59),
                        .Slide_data_60(in_data_to_next_pe_1_60),.Slide_data_61(in_data_to_next_pe_1_61),
                        .Slide_data_62(in_data_to_next_pe_1_62),.Slide_data_63(in_data_to_next_pe_1_63),
                        .result(o_1),
                        .in_data_to_next_pe_0(in_data_to_next_pe_2_0), .in_data_to_next_pe_1(in_data_to_next_pe_2_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_2_2), .in_data_to_next_pe_3(in_data_to_next_pe_2_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_2_4), .in_data_to_next_pe_5(in_data_to_next_pe_2_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_2_6), .in_data_to_next_pe_7(in_data_to_next_pe_2_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_2_8), .in_data_to_next_pe_9(in_data_to_next_pe_2_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_2_10), .in_data_to_next_pe_11(in_data_to_next_pe_2_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_2_12), .in_data_to_next_pe_13(in_data_to_next_pe_2_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_2_14), .in_data_to_next_pe_15(in_data_to_next_pe_2_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_2_16), .in_data_to_next_pe_17(in_data_to_next_pe_2_17), 
                        .in_data_to_next_pe_18(in_data_to_next_pe_2_18), .in_data_to_next_pe_19(in_data_to_next_pe_2_19), 
                        .in_data_to_next_pe_20(in_data_to_next_pe_2_20), .in_data_to_next_pe_21(in_data_to_next_pe_2_21), 
                        .in_data_to_next_pe_22(in_data_to_next_pe_2_22), .in_data_to_next_pe_23(in_data_to_next_pe_2_23), 
                        .in_data_to_next_pe_24(in_data_to_next_pe_2_24), .in_data_to_next_pe_25(in_data_to_next_pe_2_25), 
                        .in_data_to_next_pe_26(in_data_to_next_pe_2_26), .in_data_to_next_pe_27(in_data_to_next_pe_2_27), 
                        .in_data_to_next_pe_28(in_data_to_next_pe_2_28), .in_data_to_next_pe_29(in_data_to_next_pe_2_29), 
                        .in_data_to_next_pe_30(in_data_to_next_pe_2_30), .in_data_to_next_pe_31(in_data_to_next_pe_2_31),
                        .in_data_to_next_pe_32(in_data_to_next_pe_2_32), .in_data_to_next_pe_33(in_data_to_next_pe_2_33), 
                        .in_data_to_next_pe_34(in_data_to_next_pe_2_34), .in_data_to_next_pe_35(in_data_to_next_pe_2_35), 
                        .in_data_to_next_pe_36(in_data_to_next_pe_2_36), .in_data_to_next_pe_37(in_data_to_next_pe_2_37), 
                        .in_data_to_next_pe_38(in_data_to_next_pe_2_38), .in_data_to_next_pe_39(in_data_to_next_pe_2_39), 
                        .in_data_to_next_pe_40(in_data_to_next_pe_2_40), .in_data_to_next_pe_41(in_data_to_next_pe_2_41), 
                        .in_data_to_next_pe_42(in_data_to_next_pe_2_42), .in_data_to_next_pe_43(in_data_to_next_pe_2_43), 
                        .in_data_to_next_pe_44(in_data_to_next_pe_2_44), .in_data_to_next_pe_45(in_data_to_next_pe_2_45), 
                        .in_data_to_next_pe_46(in_data_to_next_pe_2_46), .in_data_to_next_pe_47(in_data_to_next_pe_2_47), 
                        .in_data_to_next_pe_48(in_data_to_next_pe_2_48), .in_data_to_next_pe_49(in_data_to_next_pe_2_49), 
                        .in_data_to_next_pe_50(in_data_to_next_pe_2_50), .in_data_to_next_pe_51(in_data_to_next_pe_2_51), 
                        .in_data_to_next_pe_52(in_data_to_next_pe_2_52), .in_data_to_next_pe_53(in_data_to_next_pe_2_53), 
                        .in_data_to_next_pe_54(in_data_to_next_pe_2_54), .in_data_to_next_pe_55(in_data_to_next_pe_2_55), 
                        .in_data_to_next_pe_56(in_data_to_next_pe_2_56), .in_data_to_next_pe_57(in_data_to_next_pe_2_57), 
                        .in_data_to_next_pe_58(in_data_to_next_pe_2_58), .in_data_to_next_pe_59(in_data_to_next_pe_2_59), 
                        .in_data_to_next_pe_60(in_data_to_next_pe_2_60), .in_data_to_next_pe_61(in_data_to_next_pe_2_61), 
                        .in_data_to_next_pe_62(in_data_to_next_pe_2_62), .in_data_to_next_pe_63(in_data_to_next_pe_2_63), 
                        .next_row_en(row_2_en)  
);

        PE_Row_B6   PE_R2_B6(   .clk(clk), .rst_n(rst_n), .new_weight_val(new_weight_val[2]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3), 
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11), 
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19), 
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23), 
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27), 
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .w_32(w_32), .w_33(w_33), .w_34(w_34), .w_35(w_35), 
                        .w_36(w_36), .w_37(w_37), .w_38(w_38), .w_39(w_39), 
                        .w_40(w_40), .w_41(w_41), .w_42(w_42), .w_43(w_43), 
                        .w_44(w_44), .w_45(w_45), .w_46(w_46), .w_47(w_47), 
                        .w_48(w_48), .w_49(w_49), .w_50(w_50), .w_51(w_51), 
                        .w_52(w_52), .w_53(w_53), .w_54(w_54), .w_55(w_55), 
                        .w_56(w_56), .w_57(w_57), .w_58(w_58), .w_59(w_59), 
                        .w_60(w_60), .w_61(w_61), .w_62(w_62), .w_63(w_63),  
                        .Slide_data_0(in_data_to_next_pe_2_0),.Slide_data_1(in_data_to_next_pe_2_1),
                        .Slide_data_2(in_data_to_next_pe_2_2),.Slide_data_3(in_data_to_next_pe_2_3),
                        .Slide_data_4(in_data_to_next_pe_2_4),.Slide_data_5(in_data_to_next_pe_2_5),
                        .Slide_data_6(in_data_to_next_pe_2_6),.Slide_data_7(in_data_to_next_pe_2_7),
                        .Slide_data_8(in_data_to_next_pe_2_8),.Slide_data_9(in_data_to_next_pe_2_9),
                        .Slide_data_10(in_data_to_next_pe_2_10),.Slide_data_11(in_data_to_next_pe_2_11),
                        .Slide_data_12(in_data_to_next_pe_2_12),.Slide_data_13(in_data_to_next_pe_2_13),
                        .Slide_data_14(in_data_to_next_pe_2_14),.Slide_data_15(in_data_to_next_pe_2_15),
                        .Slide_data_16(in_data_to_next_pe_2_16),.Slide_data_17(in_data_to_next_pe_2_17),
                        .Slide_data_18(in_data_to_next_pe_2_18),.Slide_data_19(in_data_to_next_pe_2_19),
                        .Slide_data_20(in_data_to_next_pe_2_20),.Slide_data_21(in_data_to_next_pe_2_21),
                        .Slide_data_22(in_data_to_next_pe_2_22),.Slide_data_23(in_data_to_next_pe_2_23),
                        .Slide_data_24(in_data_to_next_pe_2_24),.Slide_data_25(in_data_to_next_pe_2_25),
                        .Slide_data_26(in_data_to_next_pe_2_26),.Slide_data_27(in_data_to_next_pe_2_27),
                        .Slide_data_28(in_data_to_next_pe_2_28),.Slide_data_29(in_data_to_next_pe_2_29),
                        .Slide_data_30(in_data_to_next_pe_2_30),.Slide_data_31(in_data_to_next_pe_2_31),
                        .Slide_data_32(in_data_to_next_pe_2_32),.Slide_data_33(in_data_to_next_pe_2_33),
                        .Slide_data_34(in_data_to_next_pe_2_34),.Slide_data_35(in_data_to_next_pe_2_35),
                        .Slide_data_36(in_data_to_next_pe_2_36),.Slide_data_37(in_data_to_next_pe_2_37),
                        .Slide_data_38(in_data_to_next_pe_2_38),.Slide_data_39(in_data_to_next_pe_2_39),
                        .Slide_data_40(in_data_to_next_pe_2_40),.Slide_data_41(in_data_to_next_pe_2_41),
                        .Slide_data_42(in_data_to_next_pe_2_42),.Slide_data_43(in_data_to_next_pe_2_43),
                        .Slide_data_44(in_data_to_next_pe_2_44),.Slide_data_45(in_data_to_next_pe_2_45),
                        .Slide_data_46(in_data_to_next_pe_2_46),.Slide_data_47(in_data_to_next_pe_2_47),
                        .Slide_data_48(in_data_to_next_pe_2_48),.Slide_data_49(in_data_to_next_pe_2_49),
                        .Slide_data_50(in_data_to_next_pe_2_50),.Slide_data_51(in_data_to_next_pe_2_51),
                        .Slide_data_52(in_data_to_next_pe_2_52),.Slide_data_53(in_data_to_next_pe_2_53),
                        .Slide_data_54(in_data_to_next_pe_2_54),.Slide_data_55(in_data_to_next_pe_2_55),
                        .Slide_data_56(in_data_to_next_pe_2_56),.Slide_data_57(in_data_to_next_pe_2_57),
                        .Slide_data_58(in_data_to_next_pe_2_58),.Slide_data_59(in_data_to_next_pe_2_59),
                        .Slide_data_60(in_data_to_next_pe_2_60),.Slide_data_61(in_data_to_next_pe_2_61),
                        .Slide_data_62(in_data_to_next_pe_2_62),.Slide_data_63(in_data_to_next_pe_2_63),
                        .result(o_2),
                        .in_data_to_next_pe_0(in_data_to_next_pe_3_0), .in_data_to_next_pe_1(in_data_to_next_pe_3_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_3_2), .in_data_to_next_pe_3(in_data_to_next_pe_3_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_3_4), .in_data_to_next_pe_5(in_data_to_next_pe_3_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_3_6), .in_data_to_next_pe_7(in_data_to_next_pe_3_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_3_8), .in_data_to_next_pe_9(in_data_to_next_pe_3_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_3_10), .in_data_to_next_pe_11(in_data_to_next_pe_3_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_3_12), .in_data_to_next_pe_13(in_data_to_next_pe_3_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_3_14), .in_data_to_next_pe_15(in_data_to_next_pe_3_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_3_16), .in_data_to_next_pe_17(in_data_to_next_pe_3_17), 
                        .in_data_to_next_pe_18(in_data_to_next_pe_3_18), .in_data_to_next_pe_19(in_data_to_next_pe_3_19), 
                        .in_data_to_next_pe_20(in_data_to_next_pe_3_20), .in_data_to_next_pe_21(in_data_to_next_pe_3_21), 
                        .in_data_to_next_pe_22(in_data_to_next_pe_3_22), .in_data_to_next_pe_23(in_data_to_next_pe_3_23), 
                        .in_data_to_next_pe_24(in_data_to_next_pe_3_24), .in_data_to_next_pe_25(in_data_to_next_pe_3_25), 
                        .in_data_to_next_pe_26(in_data_to_next_pe_3_26), .in_data_to_next_pe_27(in_data_to_next_pe_3_27), 
                        .in_data_to_next_pe_28(in_data_to_next_pe_3_28), .in_data_to_next_pe_29(in_data_to_next_pe_3_29), 
                        .in_data_to_next_pe_30(in_data_to_next_pe_3_30), .in_data_to_next_pe_31(in_data_to_next_pe_3_31),
                        .in_data_to_next_pe_32(in_data_to_next_pe_3_32), .in_data_to_next_pe_33(in_data_to_next_pe_3_33), 
                        .in_data_to_next_pe_34(in_data_to_next_pe_3_34), .in_data_to_next_pe_35(in_data_to_next_pe_3_35), 
                        .in_data_to_next_pe_36(in_data_to_next_pe_3_36), .in_data_to_next_pe_37(in_data_to_next_pe_3_37), 
                        .in_data_to_next_pe_38(in_data_to_next_pe_3_38), .in_data_to_next_pe_39(in_data_to_next_pe_3_39), 
                        .in_data_to_next_pe_40(in_data_to_next_pe_3_40), .in_data_to_next_pe_41(in_data_to_next_pe_3_41), 
                        .in_data_to_next_pe_42(in_data_to_next_pe_3_42), .in_data_to_next_pe_43(in_data_to_next_pe_3_43), 
                        .in_data_to_next_pe_44(in_data_to_next_pe_3_44), .in_data_to_next_pe_45(in_data_to_next_pe_3_45), 
                        .in_data_to_next_pe_46(in_data_to_next_pe_3_46), .in_data_to_next_pe_47(in_data_to_next_pe_3_47), 
                        .in_data_to_next_pe_48(in_data_to_next_pe_3_48), .in_data_to_next_pe_49(in_data_to_next_pe_3_49), 
                        .in_data_to_next_pe_50(in_data_to_next_pe_3_50), .in_data_to_next_pe_51(in_data_to_next_pe_3_51), 
                        .in_data_to_next_pe_52(in_data_to_next_pe_3_52), .in_data_to_next_pe_53(in_data_to_next_pe_3_53), 
                        .in_data_to_next_pe_54(in_data_to_next_pe_3_54), .in_data_to_next_pe_55(in_data_to_next_pe_3_55), 
                        .in_data_to_next_pe_56(in_data_to_next_pe_3_56), .in_data_to_next_pe_57(in_data_to_next_pe_3_57), 
                        .in_data_to_next_pe_58(in_data_to_next_pe_3_58), .in_data_to_next_pe_59(in_data_to_next_pe_3_59), 
                        .in_data_to_next_pe_60(in_data_to_next_pe_3_60), .in_data_to_next_pe_61(in_data_to_next_pe_3_61), 
                        .in_data_to_next_pe_62(in_data_to_next_pe_3_62), .in_data_to_next_pe_63(in_data_to_next_pe_3_63), 
                        .next_row_en(row_3_en)  
); 
        
        PE_Row_B6   PE_R3_B6(   .clk(clk), .rst_n(rst_n), .new_weight_val(new_weight_val[3]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3), 
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11), 
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19), 
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23), 
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27), 
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .w_32(w_32), .w_33(w_33), .w_34(w_34), .w_35(w_35), 
                        .w_36(w_36), .w_37(w_37), .w_38(w_38), .w_39(w_39), 
                        .w_40(w_40), .w_41(w_41), .w_42(w_42), .w_43(w_43), 
                        .w_44(w_44), .w_45(w_45), .w_46(w_46), .w_47(w_47), 
                        .w_48(w_48), .w_49(w_49), .w_50(w_50), .w_51(w_51), 
                        .w_52(w_52), .w_53(w_53), .w_54(w_54), .w_55(w_55), 
                        .w_56(w_56), .w_57(w_57), .w_58(w_58), .w_59(w_59), 
                        .w_60(w_60), .w_61(w_61), .w_62(w_62), .w_63(w_63),  
                        .Slide_data_0(in_data_to_next_pe_3_0),.Slide_data_1(in_data_to_next_pe_3_1),
                        .Slide_data_2(in_data_to_next_pe_3_2),.Slide_data_3(in_data_to_next_pe_3_3),
                        .Slide_data_4(in_data_to_next_pe_3_4),.Slide_data_5(in_data_to_next_pe_3_5),
                        .Slide_data_6(in_data_to_next_pe_3_6),.Slide_data_7(in_data_to_next_pe_3_7),
                        .Slide_data_8(in_data_to_next_pe_3_8),.Slide_data_9(in_data_to_next_pe_3_9),
                        .Slide_data_10(in_data_to_next_pe_3_10),.Slide_data_11(in_data_to_next_pe_3_11),
                        .Slide_data_12(in_data_to_next_pe_3_12),.Slide_data_13(in_data_to_next_pe_3_13),
                        .Slide_data_14(in_data_to_next_pe_3_14),.Slide_data_15(in_data_to_next_pe_3_15),
                        .Slide_data_16(in_data_to_next_pe_3_16),.Slide_data_17(in_data_to_next_pe_3_17),
                        .Slide_data_18(in_data_to_next_pe_3_18),.Slide_data_19(in_data_to_next_pe_3_19),
                        .Slide_data_20(in_data_to_next_pe_3_20),.Slide_data_21(in_data_to_next_pe_3_21),
                        .Slide_data_22(in_data_to_next_pe_3_22),.Slide_data_23(in_data_to_next_pe_3_23),
                        .Slide_data_24(in_data_to_next_pe_3_24),.Slide_data_25(in_data_to_next_pe_3_25),
                        .Slide_data_26(in_data_to_next_pe_3_26),.Slide_data_27(in_data_to_next_pe_3_27),
                        .Slide_data_28(in_data_to_next_pe_3_28),.Slide_data_29(in_data_to_next_pe_3_29),
                        .Slide_data_30(in_data_to_next_pe_3_30),.Slide_data_31(in_data_to_next_pe_3_31),
                        .Slide_data_32(in_data_to_next_pe_3_32),.Slide_data_33(in_data_to_next_pe_3_33),
                        .Slide_data_34(in_data_to_next_pe_3_34),.Slide_data_35(in_data_to_next_pe_3_35),
                        .Slide_data_36(in_data_to_next_pe_3_36),.Slide_data_37(in_data_to_next_pe_3_37),
                        .Slide_data_38(in_data_to_next_pe_3_38),.Slide_data_39(in_data_to_next_pe_3_39),
                        .Slide_data_40(in_data_to_next_pe_3_40),.Slide_data_41(in_data_to_next_pe_3_41),
                        .Slide_data_42(in_data_to_next_pe_3_42),.Slide_data_43(in_data_to_next_pe_3_43),
                        .Slide_data_44(in_data_to_next_pe_3_44),.Slide_data_45(in_data_to_next_pe_3_45),
                        .Slide_data_46(in_data_to_next_pe_3_46),.Slide_data_47(in_data_to_next_pe_3_47),
                        .Slide_data_48(in_data_to_next_pe_3_48),.Slide_data_49(in_data_to_next_pe_3_49),
                        .Slide_data_50(in_data_to_next_pe_3_50),.Slide_data_51(in_data_to_next_pe_3_51),
                        .Slide_data_52(in_data_to_next_pe_3_52),.Slide_data_53(in_data_to_next_pe_3_53),
                        .Slide_data_54(in_data_to_next_pe_3_54),.Slide_data_55(in_data_to_next_pe_3_55),
                        .Slide_data_56(in_data_to_next_pe_3_56),.Slide_data_57(in_data_to_next_pe_3_57),
                        .Slide_data_58(in_data_to_next_pe_3_58),.Slide_data_59(in_data_to_next_pe_3_59),
                        .Slide_data_60(in_data_to_next_pe_3_60),.Slide_data_61(in_data_to_next_pe_3_61),
                        .Slide_data_62(in_data_to_next_pe_3_62),.Slide_data_63(in_data_to_next_pe_3_63),
                        .result(o_3),
                        .in_data_to_next_pe_0(in_data_to_next_pe_4_0), .in_data_to_next_pe_1(in_data_to_next_pe_4_1),
                        .in_data_to_next_pe_2(in_data_to_next_pe_4_2), .in_data_to_next_pe_3(in_data_to_next_pe_4_3),
                        .in_data_to_next_pe_4(in_data_to_next_pe_4_4), .in_data_to_next_pe_5(in_data_to_next_pe_4_5),
                        .in_data_to_next_pe_6(in_data_to_next_pe_4_6), .in_data_to_next_pe_7(in_data_to_next_pe_4_7),
                        .in_data_to_next_pe_8(in_data_to_next_pe_4_8), .in_data_to_next_pe_9(in_data_to_next_pe_4_9),
                        .in_data_to_next_pe_10(in_data_to_next_pe_4_10), .in_data_to_next_pe_11(in_data_to_next_pe_4_11),
                        .in_data_to_next_pe_12(in_data_to_next_pe_4_12), .in_data_to_next_pe_13(in_data_to_next_pe_4_13),
                        .in_data_to_next_pe_14(in_data_to_next_pe_4_14), .in_data_to_next_pe_15(in_data_to_next_pe_4_15),
                        .in_data_to_next_pe_16(in_data_to_next_pe_4_16), .in_data_to_next_pe_17(in_data_to_next_pe_4_17), 
                        .in_data_to_next_pe_18(in_data_to_next_pe_4_18), .in_data_to_next_pe_19(in_data_to_next_pe_4_19), 
                        .in_data_to_next_pe_20(in_data_to_next_pe_4_20), .in_data_to_next_pe_21(in_data_to_next_pe_4_21), 
                        .in_data_to_next_pe_22(in_data_to_next_pe_4_22), .in_data_to_next_pe_23(in_data_to_next_pe_4_23), 
                        .in_data_to_next_pe_24(in_data_to_next_pe_4_24), .in_data_to_next_pe_25(in_data_to_next_pe_4_25), 
                        .in_data_to_next_pe_26(in_data_to_next_pe_4_26), .in_data_to_next_pe_27(in_data_to_next_pe_4_27), 
                        .in_data_to_next_pe_28(in_data_to_next_pe_4_28), .in_data_to_next_pe_29(in_data_to_next_pe_4_29), 
                        .in_data_to_next_pe_30(in_data_to_next_pe_4_30), .in_data_to_next_pe_31(in_data_to_next_pe_4_31),
                        .in_data_to_next_pe_32(in_data_to_next_pe_4_32), .in_data_to_next_pe_33(in_data_to_next_pe_4_33), 
                        .in_data_to_next_pe_34(in_data_to_next_pe_4_34), .in_data_to_next_pe_35(in_data_to_next_pe_4_35), 
                        .in_data_to_next_pe_36(in_data_to_next_pe_4_36), .in_data_to_next_pe_37(in_data_to_next_pe_4_37), 
                        .in_data_to_next_pe_38(in_data_to_next_pe_4_38), .in_data_to_next_pe_39(in_data_to_next_pe_4_39), 
                        .in_data_to_next_pe_40(in_data_to_next_pe_4_40), .in_data_to_next_pe_41(in_data_to_next_pe_4_41), 
                        .in_data_to_next_pe_42(in_data_to_next_pe_4_42), .in_data_to_next_pe_43(in_data_to_next_pe_4_43), 
                        .in_data_to_next_pe_44(in_data_to_next_pe_4_44), .in_data_to_next_pe_45(in_data_to_next_pe_4_45), 
                        .in_data_to_next_pe_46(in_data_to_next_pe_4_46), .in_data_to_next_pe_47(in_data_to_next_pe_4_47), 
                        .in_data_to_next_pe_48(in_data_to_next_pe_4_48), .in_data_to_next_pe_49(in_data_to_next_pe_4_49), 
                        .in_data_to_next_pe_50(in_data_to_next_pe_4_50), .in_data_to_next_pe_51(in_data_to_next_pe_4_51), 
                        .in_data_to_next_pe_52(in_data_to_next_pe_4_52), .in_data_to_next_pe_53(in_data_to_next_pe_4_53), 
                        .in_data_to_next_pe_54(in_data_to_next_pe_4_54), .in_data_to_next_pe_55(in_data_to_next_pe_4_55), 
                        .in_data_to_next_pe_56(in_data_to_next_pe_4_56), .in_data_to_next_pe_57(in_data_to_next_pe_4_57), 
                        .in_data_to_next_pe_58(in_data_to_next_pe_4_58), .in_data_to_next_pe_59(in_data_to_next_pe_4_59), 
                        .in_data_to_next_pe_60(in_data_to_next_pe_4_60), .in_data_to_next_pe_61(in_data_to_next_pe_4_61), 
                        .in_data_to_next_pe_62(in_data_to_next_pe_4_62), .in_data_to_next_pe_63(in_data_to_next_pe_4_63), 
                        .next_row_en(row_4_en)  
); 
        
        PE_Row_B6   PE_R4_B6(   .clk(clk), .rst_n(rst_n), .new_weight_val(new_weight_val[4]),
                        .w_0(w_0), .w_1(w_1), .w_2(w_2), .w_3(w_3), 
                        .w_4(w_4), .w_5(w_5), .w_6(w_6), .w_7(w_7),
                        .w_8(w_8), .w_9(w_9), .w_10(w_10), .w_11(w_11), 
                        .w_12(w_12), .w_13(w_13), .w_14(w_14), .w_15(w_15),
                        .w_16(w_16), .w_17(w_17), .w_18(w_18), .w_19(w_19), 
                        .w_20(w_20), .w_21(w_21), .w_22(w_22), .w_23(w_23), 
                        .w_24(w_24), .w_25(w_25), .w_26(w_26), .w_27(w_27), 
                        .w_28(w_28), .w_29(w_29), .w_30(w_30), .w_31(w_31),
                        .w_32(w_32), .w_33(w_33), .w_34(w_34), .w_35(w_35), 
                        .w_36(w_36), .w_37(w_37), .w_38(w_38), .w_39(w_39), 
                        .w_40(w_40), .w_41(w_41), .w_42(w_42), .w_43(w_43), 
                        .w_44(w_44), .w_45(w_45), .w_46(w_46), .w_47(w_47), 
                        .w_48(w_48), .w_49(w_49), .w_50(w_50), .w_51(w_51), 
                        .w_52(w_52), .w_53(w_53), .w_54(w_54), .w_55(w_55), 
                        .w_56(w_56), .w_57(w_57), .w_58(w_58), .w_59(w_59), 
                        .w_60(w_60), .w_61(w_61), .w_62(w_62), .w_63(w_63),  
                        .Slide_data_0(in_data_to_next_pe_4_0),.Slide_data_1(in_data_to_next_pe_4_1),
                        .Slide_data_2(in_data_to_next_pe_4_2),.Slide_data_3(in_data_to_next_pe_4_3),
                        .Slide_data_4(in_data_to_next_pe_4_4),.Slide_data_5(in_data_to_next_pe_4_5),
                        .Slide_data_6(in_data_to_next_pe_4_6),.Slide_data_7(in_data_to_next_pe_4_7),
                        .Slide_data_8(in_data_to_next_pe_4_8),.Slide_data_9(in_data_to_next_pe_4_9),
                        .Slide_data_10(in_data_to_next_pe_4_10),.Slide_data_11(in_data_to_next_pe_4_11),
                        .Slide_data_12(in_data_to_next_pe_4_12),.Slide_data_13(in_data_to_next_pe_4_13),
                        .Slide_data_14(in_data_to_next_pe_4_14),.Slide_data_15(in_data_to_next_pe_4_15),
                        .Slide_data_16(in_data_to_next_pe_4_16),.Slide_data_17(in_data_to_next_pe_4_17),
                        .Slide_data_18(in_data_to_next_pe_4_18),.Slide_data_19(in_data_to_next_pe_4_19),
                        .Slide_data_20(in_data_to_next_pe_4_20),.Slide_data_21(in_data_to_next_pe_4_21),
                        .Slide_data_22(in_data_to_next_pe_4_22),.Slide_data_23(in_data_to_next_pe_4_23),
                        .Slide_data_24(in_data_to_next_pe_4_24),.Slide_data_25(in_data_to_next_pe_4_25),
                        .Slide_data_26(in_data_to_next_pe_4_26),.Slide_data_27(in_data_to_next_pe_4_27),
                        .Slide_data_28(in_data_to_next_pe_4_28),.Slide_data_29(in_data_to_next_pe_4_29),
                        .Slide_data_30(in_data_to_next_pe_4_30),.Slide_data_31(in_data_to_next_pe_4_31),
                        .Slide_data_32(in_data_to_next_pe_4_32),.Slide_data_33(in_data_to_next_pe_4_33),
                        .Slide_data_34(in_data_to_next_pe_4_34),.Slide_data_35(in_data_to_next_pe_4_35),
                        .Slide_data_36(in_data_to_next_pe_4_36),.Slide_data_37(in_data_to_next_pe_4_37),
                        .Slide_data_38(in_data_to_next_pe_4_38),.Slide_data_39(in_data_to_next_pe_4_39),
                        .Slide_data_40(in_data_to_next_pe_4_40),.Slide_data_41(in_data_to_next_pe_4_41),
                        .Slide_data_42(in_data_to_next_pe_4_42),.Slide_data_43(in_data_to_next_pe_4_43),
                        .Slide_data_44(in_data_to_next_pe_4_44),.Slide_data_45(in_data_to_next_pe_4_45),
                        .Slide_data_46(in_data_to_next_pe_4_46),.Slide_data_47(in_data_to_next_pe_4_47),
                        .Slide_data_48(in_data_to_next_pe_4_48),.Slide_data_49(in_data_to_next_pe_4_49),
                        .Slide_data_50(in_data_to_next_pe_4_50),.Slide_data_51(in_data_to_next_pe_4_51),
                        .Slide_data_52(in_data_to_next_pe_4_52),.Slide_data_53(in_data_to_next_pe_4_53),
                        .Slide_data_54(in_data_to_next_pe_4_54),.Slide_data_55(in_data_to_next_pe_4_55),
                        .Slide_data_56(in_data_to_next_pe_4_56),.Slide_data_57(in_data_to_next_pe_4_57),
                        .Slide_data_58(in_data_to_next_pe_4_58),.Slide_data_59(in_data_to_next_pe_4_59),
                        .Slide_data_60(in_data_to_next_pe_4_60),.Slide_data_61(in_data_to_next_pe_4_61),
                        .Slide_data_62(in_data_to_next_pe_4_62),.Slide_data_63(in_data_to_next_pe_4_63),
                        .result(o_4)
); 
        
   
endmodule
